SR    
  h                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           Tue May  6 12:24:51 2025   sboardse   (gs674-boardmba-198120187032.ndc.nasa.gov     �              arm64      darwin     9.1.0       ��           OUTS2         4      נ   z                 z                        	          !                                                                        	       0          8          @          H          P          X          `   	       p          x          �   	       �   	       �   	       �   	       �   	      �   	              0   	      @         H         P        �        �   	        	     0   	     P   	     �   	      DABS   DDXX   ICON   IERR   IRK    ITER   FRQ    FCP    WC1    C      VREF   CINDEX     WNA    X      Z      P      D      DX     DZ     DP     EFL    BFL    VG     XX1    PP1    ZZ1    AMU    DN0    DNS    VS     JS     XES    EDIE         0                                                  0                                                                                                    0                                                  0                                                  `                                                                                                                                                     @   $                                              �                                            @zJ{��-=o�nq              @� ��ǫX>Q�{7:�@���	| f@��8�%wA��xt   @�8`uR�N@� 9�@V|�����@��b傖=��*rX�!>�s��S0?�Į,�<��zJ     ��Xx  B�����A��d�~�U-?�-����_8j��Q��Ɖ?���9px�?��3�La        =S����?����3}8?
�~ݯ�ٽ��`��d���K+�@:�sX���j?V�L�~��=�w��w��=k���=�?�⧲@�@`W�,0^@cA�+�@��b�j�=��)ui>�?�Į,�<�>�s��S0?�      @/��[W>�                                A�e��@  BL+��  BL��                           >����A@����{�>��xc� A�y�*K>�r�M��jA+|�s                                                =�5�>J1@Lv29e@pH�ƪ��W��
�>f��	��?7���`$=�l���?�H@�ڪ�b�]gu�=0���
J>e��>���ל����r�jsG?��挕]�5 �T�3=�Wȍ�q>LP��ہ��&��                                                                                                                                                ;��f+B>:�ۅ��p> }�Ԣ�#�����ت<�&X�
2=T	{��_<U���#>R8I,�r�اN�?e�;��c��<z��$�C=n����GG<tx�Xi7�X���s�>����˟y�p��a.��ĩ��0�>\	$�>�i                                                                                                                                                �I�4O��>��Hu�ȾIm~V��15�-�%���m���>�������I��4��H>�=�^�K>x���%:�>��f�����F�0����v���a��Pk@>"��O�l]��xr
��k�V������w���4>�: �q�h�a�����>"��0拏>0�A��>I�)��}�a���_80>6�� @@&\��  >,��W  �j�jL����ƾQ���6�I���y�qn@!��  >1pf9�  ?c9��YE�?��%*���P];����<?ͯ�                                                                                                                                                                                                                                                                                                �fs�wT� ><���� �k'�YS}/���ỉ�̾ȴ�%�˾�6�2��f�`��  >?���U� ?c9��Yek?����� �P�z����<?�V�@x�1��� �DJ��r�>k#�-v�l@���;3>�e��" �>���c��@y�8a{Z�H�����s:*E��B���,�A`��(5�?��2��w־
����2�>0Yb��0���q��R�&>I�P�V�ȴ�1�����c�7}�쾘5�,�
>3Ls<���+T��e�w?��]	)M����
��X��\R(�d��������=�όpV������h��g>,[�9����<'��ξ�6����lNB)�>�(N��?c9���-�?�ߺ;PR@]�^�L0>9��R�M}BG$Iѷ�I<��8O��$              @���<;j�>��
e��@���	| f@��8�%wA��xt   @�8`uR�NAB���N�@V|�����@����>>� x�×?xX�_���@>���Ɩ�FhD�$ �,�5��]E.�`$��C��\X�D�g� b����P$��SD�ɤʟ{CP�}�љ�?���3�k�        ���j�ed�>��R\�G?L�L�g⼽��+'}�?<ݠ:�ؿ�q�l �K?�JyΟ>T
�;1𽀓��jr?!�5^��sv"̋�������8|@����t>>��+#@>���Ɩ?xX�_���?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?���x��#A^m�1��@0 8X��P0�2|�@1z�q�)�AIO�Lg'�                                                >�o�^�z@��A��N��
h�V�>k����>���b?�+G=Ӓ>��#s
�����Ug�ҳ�9��>�X��>����4?�_�XcB���4;�n�r?��j�Q�4K�f���x�h`��?$8A<Q�.�%}�                                                                                                                                                 <��U��>$�MʞH�)%��<��@�7+<�Y�-��=�Cc��<���-2XR�4^{������|��~��s�i=6$�,.��>x�o<MoA�����'Hv>��T�U�=	�ۋķ�������>�|]?���                                                                                                                                                �3@ޥ��@>���N�>�{J@�WB@�� .Z�����A�~?#�E^�^�V�^A�,>�FF<�*��;��*��=�j�T��V2��?U-)��@$�/��AP?���	E{����[goj@"��:�"�(;�+شC?D�Q}s��_ٿs�\>�Qq��]? �:��;�?�x�����_�OUf�`U���i�@%�e�  >����� ��gQ��iv���{�5*?�A|'���w�R��.|n��	�m�T���`��Ĭ�������@�Ӫ�[���Mt�H�'c�K8xD�                                                                                                                                                                                                                                                                                                @�b�  ?A�6 ��ҁ�K�����e���+� ҿ���@9/��	�#�T �`����~ȿ���)�@�Ӻ�^��Mu(f���Kx�~�	@��S �>�?�aY"�=i��ܖ����@Ƃ���n����ވ֟���^e���A�7�S�?�7�m��@.@UH=MZ�ULA7�A^7J-O}@�!�/mW$@7�\W�?&��,��b���?�t�kC�.7!2)s�Q"r����Z��#�����Vu��{U��@����
��'"�T�A�}l�()�@�G#���? P8�.������,@�HN�̕��J�w��n$?W,������	V�o�n��)/��n��!"E@�6S�B�A
��E?@�WTs�*@n2��jd=eM7[>              @����	��>S�5�N�@���	| f@��8�%wA��xt   @�8`uR�N@�(έ�B@V|�����@�v|ȏ=���gT��>�PU����?��y�A�/@n2     ���_m�  B���
A���Q.*�S��%g���[��
$�L�[!�C}�����C��?��s�5=        =S_�h�l?���
�F�?/s�ȼ ��QyKࡼɷ�?J�������?V�2�ε�=�{�X<�=lǮ�w��?��Z(n�@_��O%g@d�Ɨ���@�v|�&=���i�j?��y�A�/>�PU����?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�L�I�@�ֲ"{�>�AT���AX:�)h>�-E�zS
A㺐�m�                                                =�4���@���+:A@��l),s�Ѷ�\/��>e��&�׃?8�l��#=�D��},�?���	c2*�`�ۇ[��=/�qq�->�C�KF>���yP4����~w�%?����,�5 E�ŋ6=��_	\�>MS�٦Nؿ�N��                                                                                                                                                ;�A����>9NY���
>7s�訳�����Z<�Q�?��=T�	�=�<n��K��>Q�랗g����� �Y�;��sj���<y����0|=o��{�<
H�dU��W�n��G�>���2ϼrK@�]���pcs��J>]<��㘌                                                                                                                                                �G����%�>Emk%��VY͞�.J�E�ɾÎ�K%�>���3��G�58��d>D�Y5��>u�sͿ�>�1X�8�E'�������f}���`4��l>#K�T57����2+#p�νs�������>�gj�rı�`4���>#K�'}_>.��Y�>G7�g[��`2fG���>
c�!��@&\�  >,ͯ�� �l����������8�?�ӧ���� Op@!��B�  >1��(�  ?b��2?�	'��M�==�ʿ����)�                                                                                                                                                                                                                                                                                                �d��Q� ><�!��  �l�r�dG���vKY6<�ƞ��oi�̤u�$�d���� >@�ᠠ ?b��)���?�f��M���.�s����m�U@v�4���w�G�R���Z>mӸ=��2@��jOd$�>���eo��>��U_��@w&�*�Lq!4� ;�r�L�U$�MؤA]����?��i*R��,VĀ�G>09���]���*@����6���E �ƞ��U���D�����6~��9>35�%W�*�r��A?����տ�l(��CE�����|����gvQ��>#�#���{"���2��`������Ƣ@
�,~�̣�Sd����`N�>'o���5?b���Ǧ?�
H��7@��5�c>9��CO:�Be�N[fYf=	<��<NL              @�[�X�>��YY�#�@���	| f@��8�%wA��xt   @�8`uR�NAѫ��S�@V|�����@	������>B鳊�{?<m�s'�@!z;��iBe���$	 A������E0��A�I�C�=�D�7L��½�"wT�!U 5i�D�l�K;CqP%4�?���3��_        �4��`n�>�⎭�?L����R����~X='F�i�v�w����P�?����)0>&اM��o�@.�?��/��L�ql�h��g?����):@	�����?>B鳘��@!z;��i?<m�s'�?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?��D�p��#zgZ@Q���YAT�l{�1@R
��wxAPd(�!�P                                                >z#�9a`��qj~Yd��CF���>H"�������m���?r?����cAh>���Z
/�?���3Y濐l �ʾO��:FA>�s6f�w~?��Hݯ�$��D�@i�?�M[��&��3�����C��n�"?@��A���$�l��mf                                                                                                                                                <�'�n������hi��U�,C�<dy��U�
��EQ�:�=��W<Z=�e��>��G���U��J޼����d��<�*^��8>��O�w<R���o�Cv�>�K�{�=Y����9��^��}0>�QRs��B                                                                                                                                                ?�:�If��>��0�}�&>r��6?�������ڃ)ͨ���ıe�����A�9�4�#>�
���[��E��1���(���AuI�\޾�`�ۇ}��$��y��`?!�b+𿁾�pӠ�8@��?�NZ�"��;5?
���l�^��:��z? �Fڊ���
���N?�ޱ+er�^�^�� ��2炔��@%����  >��5��  ����19��$���r�LM`t5ͿWw!q��3��r�X��o!����	s���*�@�}�����K9��Se��f�I��                                                                                                                                                                                                                                                                                                @�Y4`  ?!�M�� ��t�|:J�����q���"�&��P�VJ뤯kx�6>U�h��nO�;��	s��c8�@�}��F�H�K:*�&�0�f�X��
@�E�J�~?��8��-�B��E�B@���CY������f��?�~A>nA#Ɠ��D�?�)Dە�5@E$d1��@�4�Z�n�A\H�}[�F@�����@�v��cc��ݧ>ʦ�_.�c?���O-��#�7�ϰ�?E0�
�)����D`A����-N�i!�1����Ma@�������6�T����}����@�6�����?(+�P�>ޢ6�R@��_�^I��4�P�y1y�X6*ף��!��:'��(��֭��TjGq@��A�#K�A��ѾI�@/�L{���@q;���=l�M�b�              @�_����>Vv��a��@���	| f@��8�%wA��xt   @�8`uR�N@�$HD�'@V|�����@	���=��狂�T>�/a�1c?����=�@q;     ?�	Z�  B�LР/�NA_��Q.�g>����fs���G�-��Q�~�+�x'?���1� D        =S����?�c2�@?�"�������&���������<��r[I�?V��A�=�����U=m�?c���?�KxmU�@_���v'�@f��fnR@	�����=����O9�?����=�>�/a�1c?�      @/��[W>�                                A�e��@  BL+��  BL��                           >��n�4i�@�Z�Dd�>̲�+V2�A�+��pQ>��p!�I%A�'gd                                                =�H�,Ґ+@~���v@ `��l�%��9^����>d����V�?9� ���/=���E�?����ϫ��]�N~�C!=-��$Ȏ>#ց>���\�RŽ��D@@�?�1����.�5 k_��s=���h�j$>N]'k��տ��FSL��                                                                                                                                                ;��3M�E�>8,��$�>�9��[��9骒d"<����;/�=U�:
I��<�}B��I>P���ށ���u�iy];�|�ă�<x��'+�#=p��}��<�<�7J��V��/��M>��4�6�˼s�'�XM��� 5WX��>^p|^�m�                                                                                                                                                �E���:V^>�LP�����v|�r�*�,�8������,)��>�n������E�U���c>���gkd>sn`+�>� ��^O��C�@�e~�P�B	�s�^y��>#�Za�0�҈���F��]{t����/nf;!>��F���.�^s��>#�Q��t>*�qW��>D߽��\�^��KRn>	��5�@&\h�  >,��� �nNm?g�J���ܤjv}�;-��ۊ��-��it@!��#  >1���o� ?a�vsd��?��e���Kv���j��+�HD                                                                                                                                                                                                                                                                                                �b���  ><��7q� �n��*PO���וFh�b����s�����6�&�c4��v@ >@�_L  ?a���u:?��n��Kw
��;��+���@u� v_�G�Dx��>ot�j�@���.�{>段�Q0�>��9�]q@uNk�� H�Le*MS/�q��goy������A[w��#?��R0\�):ɗ<�>0!^}z�I��S!0L~�6��Sb۾��������%v�㺾�s���|>3&X��ɾ)��j*��?��T��{f�(\ῃMM*E/���zT����=B���D�C�s04 �u;�A���Έ�����݆��{�:�	���2P�>>�#�0Qi?a���bJ?��A~��@����T�>:�w�WB
i�[VXV<�ؒWo�>              @�	����>�v��F�@���	| f@��8�%wA��xt   @�8`uR�NA���@V|�����@
̩u�^>;k��m�4?�S`>��@&���rO�U�@ A���Yj(�E:ƽ�;��C�G8��@����(Нr(D8��x�D���,{�Ccs��K�?���3��^        �%<:�5>x�+�;_C?L�	��S��y�K�Lt=�A��T�q�'���?�����!>�]���ݽ��DYt
?Ͼ_]&�i3��� ?��G�s��@
̩u�^>;k��9�@&���rO?�S`>��?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?�����]B�C�)��@I��s��A`�[��E�@IȖ�(�AU7�K���                                                >]����ѿ䓲'����`"*��>,X��pg���� O�?�����N�>�vi��?��2A�+F��C�G;�2|/���>\�+���?�B�+͛��:�2��^?��D/;��3"�u���s8o?32�V���#���f�                                                                                                                                                <y���}�u+I�HR��"���A<HƮ��}��qU�=��zo�=���"�>������� ��Ƽ��4e�[<���z��>-�&^*�<I}�?��v��8]
>�@|���=UF���Խ�r�[|��>�"t�ii$                                                                                                                                                @<�� >�����u>T�=8��?�,�h&�����q�O ��/b����.Ҕ�M�>�dQ!�%����2zd���G_�]�-�s+N?���b��(��)��Z���?���꾴���\��@�\2�\�"�VZw>���{4��]&^X��'>��2��g辽ߥU?�?����Z\�]�ѕ�%?��r@%+��  >�J�U�  ����b�fO��M�æ�WE$@Ĺ�\M�`�;��T�I�'E��wAٱ�@����2��I#˃���W�1��                                                                                                                                                                                                                                                                                                @4w9�  ?�(駞 ��QUyw�n��I��o���#<qCۮr�\V&��8�$󗤘��H������wB�&�C@����؟�I$��\��W�/�ͺ�@�U��W?v�⣮�K��7%��R@�66u,�C���b��b��_a�K�A.��5-p�L9��L�]�Dن&����]AZ���n��v��e�?�m^Hγ�>�G蹯�_.n�!v?������#�kJ���?$�c�'ʲ��i���|@����+@O�씂�A EVҕ����b�:�@�uMn`{�@sF%���
��G��p>���\ж@���6E���kZ��\:�o���)�^�=����x���S���r�.��Z@�<~�]ABp�֐-@,���ĂP@y��1R��=xA�o��=              @��=�fi>Y�qø�
@���	| f@��8�%wA��xt   @�8`uR�N@�4����J@V|�����@
ڌ�*=���@��>>���ˆ�?��S9�T�y��    ��Q+�`  B�m�����A	��l��C�O$ւ�f��	~��0�C�����y��T��|?���"        =T�E�-.�?�R9���?�9ek����4B#���(�dn�3����?V��Ft�=����>ȡ=oF�J"&?�+�/Ri@_R~|l�@hd�>a!@
ڌ�)��=����i�?��S9�T>���ˆ�?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�;����T@�maLLp*>�%<L:@�A�&��>��2��2�A
��(�                                                =�bF˅b?@G��t?�;Z�ޢ/���՜�3�>c���!?:�`\�=��rQ܏'?�w)m8ڿZ��g(�^=-�Gú>h�f�S�>���膥I���;�$�?�������5 �����> 8p����>OlXx�[��ޟv��                                                                                                                                                ;����%��>7%ρR>�&}�%��z���N<��<)z�=V����<��5֘>PAiwA�ͽ�Q��4Y�;���U <w�ւ��=qK�&�(<�bC<�U�wI�dL>��`�J�C�u���5��������a>_�~�":�                                                                                                                                                �C������>����n��JK���'�[�=�4������)>�b����C�i$tn>��xVB�>qX9,xЫ>��'����B7�cg�'����[�D���>#��u�����3�� ��N���_��>�P$�h�[�>��S>#��eU�`>(4�h�@�>B�X�"�[��O>�խm�@&\��  >-��� �p }�d���N����=z��ˡB��>N�u�8@!�"�0  >1Ċ� ?aZ��N�?��DO�/��I�@������߆��̳                                                                                                                                                                                                                                                                                                �an�� >=J��  �p(�\ H����L��E���E#���e�`��a�G�2� >@+i�  ?aZ���"?��F }���I��|�[��߆�K&@sq�`���G��,>p��U��<@���~0W>���O�>��H7)2�@s�����L_|DB���qZ� ��B��Lu��6AY��c8޽?��fo*nξ&Ϳ�Ѳ�>0�h�78����w��5��~����E
�����dn���\��~׊kB�>3ɜBy�)8��ΐD?��F��A���B���0���F�L�����/0��`@G��F�~�cn��?Fw4�����G�ue�0��e��$�ٰ/�C> K[��?aZ��U?��D�P�@ι/6.�>:^��uB��Hf�3=k���e;              @����q�^��ͳ��@���	| f@��8�%wA��xt   @�8`uR�NAH��h��@V|�����@�ȵ��"�sj>w�T�?� �^��@.W�7��_��> A�Hf���EI�vd,.�D�SvV���u�J@�DT��i�D�8 �
�?Í;���ڽ?���3�R�        =VBb�U~>j��_%3�?L�7�e��=�h6o��Tg��ODh�h��	9<8>�oVu��7�x�p=�ՅB
��?��}+�`)i�tp?�-f4�y@�ȵ����sj>wM�@.W�7��_?� �^��?�      @/��[W>�                                A�e��@  BL+��  BL��                           ��l:JԴ��E��Q>��y��9b
pAd��k=rM�y���z�vA[g�
dE                                                �n�p�F-V��b2h�HR���&e}��7Ѣ��	㾾!�߀R^?�y\�L�_���<"��?���N��vN;�9��>D�Jc�5����e��fI?�L1=�*�>	�-�L�?�WG�L���1������?E��W�"�]���k�P�"�d���j                                                                                                                                                ���s6Z��0C����gQA�*�T5L��Ö�ِU�y��=�6z��1|M
�">�8��޽��S���
<�����ż���6�>��RƼ�#S�F���PB$�P�>�f&�N���g�9~�=Ә"���>��4���                                                                                                                                                @�2J�@�����R̾bN�@�q�?��{̔k3���ڋw���:Rtt�e�v�Kw���E�ܻ!߾�]=��Ŀ��Լ���[�B>0�ؐv�G��'��Tq�=�e K>�-9��?��"(%�&�)�#��1�^\#�[����nX�1�r��{�����
��?�e��4%�[�_��Z��EHF�̕@$1�τ  >�3R��  ?X|L;����@���c��e��auu�|�&f���	P@tP��e�@B���3�A.��#J%�G$��1@�I���q                                                                                                                                                                                                                                                                                                @���  �<��� ?��@M���:��%-�'�57iv�a�v�y�&g��D�(@t	p�/@B��׏4A.��5Z��G%%g�Ke@�I���@�P�H1?���*�`��-D8^@@�Q,mJt@~��Ll�?�.�K�A"A7gC*o1T�>j��mB��t����*j�(ågߏ�AY���C���X��"mD��WQC��Կ���>��/ӓe�gsb����'�;��gv�9�,K����̜���@54[\���@`aH�s�AX��g�(�%����t�@�i9rGU@@f�E��?CZ�,�O��; �:Z@���}�5@��K� �]��7*���1��%Hx@a�Zz�@5\f�fA@�E͂-�qA'��nV��b�}���@�y��v�=�^�D��              @��nځ�n>\oS�� ]@���	| f@��8�%wA��xt   @�8`uR�N@�B�ZЕ�@V|�����@�{I�Ȅ=�l�&2>�ԗ0�3;?��oqto���y�    ���K!   Bѭ0��Ai4�[Xd�L���ˋ���w�L���A+Im����u��<A�M?����ȥ        =U	%� j<?�t�ˇ
?!	�]����fX/���e;CF��j��8��?V�3�1=��� =p-K��g�?�}U�e>�@_ԶOq@i�y�	L�@�{I� =�eӉ?��oqto�>�ԗ0�3;?�      @/��[W>�                                A�e��@  BL+��  BL��                           >���O�J@�y�W%�>�l	J	KAmqo{�j>׻�O_��A
��uΆ                                                =��0V�p�@P�?��?�Gd�#΁��v΍��>cC��P�?;���2�F=����d��?�Dg��ԃ�X	p��=,	m�M��>�"��>��|�%�����R�1?�W�aK�5 �e3�>V�Tp>P-���� ����                                                                                                                                                ;�c٬m>6R�3�j�>��l-�����|�<�XEv
��=WZa�B�d<	��nN�#>O����]ͽ�S��;�;�63��߷<wEV�[xy=q��/e�B<L������U8�����>�ׂ���v�@%O����r��}I�>`W��f)�                                                                                                                                                �B�+��z>\I��R� G��+y|�%��B䋏���V���>�M�Fb_�B���DQ�>[�96�>o���:>�%2��A!p1RB���Bͭ�Z=����>$Rpa��ѱ���9F��R�$�d����&А�>�*f�c���Z=}i�\>$��]>&%���>AM&����Z;FoQW�>?���q2@&\<  >-!���  �p��D6���)�<�v	�?���y�w��L�(�K�@!���D  >1����@ ?`��gn?ጣT���G�IMXj�����^��                                                                                                                                                                                                                                                                                                �`EK`�� >=/���  �p�{��.���6�bU50��O�ھͱи����`���� >@>w�A� ?`����?ጤ��6��G�daJh���˻�cl@r9K��Z�G�T�v &>qA����+@�Q��^>�m�.�>ǒ�Y0��@r��E���La]���6�p�AwO�����F�AW�eB�qU?�Y����$� ���.>0 �E�{ٽ�ow�m�5jH��T���MK���{��K�����5";�>3��ߝ��(��?)�?ጥA�%ٿ�^��ϷX���xyd����	KI�%�=o�* ��#�L�+z�ft?ZI��ޘ`��A��ݾͱ�����b���w>lJE?`����N?ጣf�K�@�Z� �>:�&�V(,B�\�J��=4q��n              @�X@n�D��qmqsbP@���	| f@��8�%wA��xt   @�8`uR�NA�U.G<z@V|�����@��8�db�؎X!��?��+��7�@5�>bZ�B�X���$S�yU�,Π>Ea��7�D�����+�.�#y��uD��rq��7D��c�7�����&]?���3���        =�"y�,ջ>VS�Y\\�?L�U�a=厪��
���x���ns�\�1��Ǜ>����2M�������>[b�3ɶ? >��ɿP��tȯ?�t�f|CS@��8�f��؎X٨�@5�>bZ�?��+��7�?�      @/��[W>�                                A�e��@  BL+��  BL��                           �)H!$�4�A֖I�v��3D���0Ah�r�v�*��4���Aa�m��+                                                ���7L��Ԧ�����W(dQO�O���?�M����l�D4?��p#�����P]+?���r�߿f�Ig^<���O��meݾ�Ȩ�H7�?�^��L>mg�R�;R?�սb���-��f>�S?�G#�ڿ���=����"=4;�z�                                                                                                                                                ��(��x��.g��
�s����g��Sì_���XPJ���=������m���N�9?E>�����ݿݜ�μ�1=2�hg�&�>$с���w��}�Qܿ��v��cD>�������� �/�s�>2�אR��>�-�� �                                                                                                                                                ?�(���`���%��bP����!�E�?�;>����9�QZ���|R�v9�?�tCv��&���8Z׾�����p���������?�晷�F��&�u^���#S(���ȿ�#�-����u�?��:]kt�0�F�_���s�KL���[K��N������0p>�%���@���*�} B�\U@�]����}1Y�@"42
x  >×���  ?y!".4P-��Vvde��q�#^�z�e�u= &�24��Da�@���A��@�!?�{AA��r�E���K�@��`�                                                                                                                                                                                                                                                                                                @�p��  ��%ς` ?x���H#��T�
�[��0��0�ڿ~�1���x�25AY^I@�K���@�!?G�\AA�����E�HWzf�@��i��@��>mjW@@�#�7q?aM��[�d@�*ă��z@����'�@ �x=IZ�ADq�^$���ɦ�����(�9���9�E�59@A]+l�Jn��!�A$�q����RkͿ]���ž�s�&;�?jQAZK��34Ã�?iv:���B�
��a�KY@�Kǽ͕@�F{�x�A !���|�=^����A��d�0�@X}��?�t��ֽ�u�;1�K@��-��@3%��T9�?oH�Pӽy�5r_�Kc�@�Eb��"@�v�R���@�o��Ca�A5����Ji��׶)Km @qn��.�t=t���lOo              @�V�t��d>`�%��@���	| f@��8�%wA��xt   @�8`uR�N@�S����@V|�����@����̮=Ə.�(k>�����*�?������qn�    ?��Ԉ  B�� �x�A�}�;�J2L��������Z�l�<�%ԧ=;�r]@w�?��0��t        =Up�!;�*?��TC��?sx软���:����ť0�� ©���?V�
2�=��G���=p�cU�1?��j���@^�*+�[@kӜ�ț@������=Ə�����?�����>�����*�?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�)'�m$@��w�v>�tX$,\A�^���>ؓ�kbsA	K� ��                                                =மB�KZ@IF^y[2?�C�B�tؽ�%=��J>b���G7�?<����j�=������b?�sK
�1�U{އ�Nd=*X3:�ڮ>`ƙt{>���a�(Ƚ�#
��h9?���Ľ�5 �#It�>������>P�=|�>%�鏫5�c�                                                                                                                                                ;�N��{ P>5s��e�Z>H�7�ǻ�e_9�'<�em��=X5W��<
�羳w%>Nw�����	�-�;���IJ<v��h?Ni=r��>��<�1����TxJ�v�n>�צPz	��x¶�D�ּ�,�I���>`�G��g$                                                                                                                                                �AYh�e�z>#���@����f#�#_˳������-��>�q�����AY-I�>##k�>lj-�@S>���-[��?��<=��aK"����X�k"	�>$L>c�Y��F�ѹ���\W�x��ʤ���>�����=��X�e��ì>$L5w��>$=D��>?xΐ�B��X~w$'^�>&��a�@&\X\  >-?�5c  �q�����k��b'F�@�A
gcu�%��]t�Z��@!�$�  >1��I�@ ?`a�	��?�KH�u��Fh5�D���zy�                                                                                                                                                                                                                                                                                                �^!�j�� >=N�9Ԁ �q�*W�@��m����G����V����OZN���^�[ɥ  >@Ub�s` ?`b�;N�?�LŁ��Fhvq��W���N�j|@p��8m%��G~�v��i>r���^,@���?oc>����-�>�Q��@qAٍ�˓�Lj�O��>�pb=*����SŊ�AVhwM�݃?��I����#/�O7?�>/���r!e����lӗ�5O���Ⱦ����:���j�����;�V��)>3�o*��(%����7?�MQ�sj���_�����i��@��8�A䌽T�������w�C$�?d��Ny������٥1���5���� ���ۗ>�6a'�u?`bf4��?�Kg�@�seWP>:�׼ˎ@}�2��=�� �+I�              @�D-}�>a��W;��@���	| f@��8�%wA��xt   @�8`uR�N@�d�Y�G@V|�����@�Ѳ��T=�K�[q)>����o �?��aڤ��@}�     ���)�  B�է[��A 8I5pc@�H���_���mނ���8��rme��oH� ׁ�?��Uq�ő        =U�a��:�?����ۀ�?��������|_�x����|���,� %��K̷?V���]�=����4=q7���
�?��9���@^}�'\�1@m��U��@�Ѳ�A�=�Ho�L?��aڤ��>����o �?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�|�rv��@騡tl�>�5���AON�~��>�b,Ț�A�W��\                                                =��9�A@WC����?�w�v�ϼ��k<f>a�[T5��?=����\�=�b L�c?֯«��ſS"�P4=([~��"
> �(8�>��ő?d���7TB3@?��\���5 �#(>����e>QI$������w6Y�؈                                                                                                                                                ;���sO>4���7|�>����V�����F�\F<~|I?Hx�=YL�}�j<ǘ���>Myj�o���<++�;���p��t<u�_�(=s-l&��<���)��S��"�^�>��� ��@�z���`߆���'C{��>a��x
��                                                                                                                                                �@&.��]�>�u�yaA����/��\�!r8�XȾ����d��>���Y�p�@%����n>��en�>i��	�>>�Ki�[b�=�Y��ӾD$)��(�V�!>$��t���������/=����W������>t�F>��N�JLK�V�+�֢>$��`�ט>"=!k�� ><���8m��V�\��->�O�q2H@&\�h  >-^%��  �r|������b�ԾB[�����n���|@!���h  >2��r  ?_ӡ�n?�^���D�]�/Q��}�ۮ�P                                                                                                                                                                                                                                                                                                �[��^T� >=n�� �r����������r?.����n\���R�H�*�\���"  >@l�)�@ ?_��HA��?�`<3��D��"D �}��m�F@o�����|�GyEH
�>r��aL@�Ǉ�u�>��� %>�	�'k�@pՖ5#�Lygl)+�o�6�9T� �fxI!�AT������?�O�n�h�!��P�aQ>/�W����� ��ƾ5S��Bx���nR�)���㢺�����߽?]>3hO!��'���SIo?�`ű�������y�}��%I�����{��=S�&!���ax~��QY?kq���������nh��Ru4���H�<3�>\~��?_�ԐON?�^̥�J@@+��|>;?LQ�3@b᜸T��=lZ�5\              @���OΦ�>d(;��@���	| f@��8�%wA��xt   @�8`uR�N@�vC[!�.@V|�����@��؛�=�8&��;>��|��?�����8@@b�    ?�wR��  B�Jp��@��I�>��F0{���(%�1�q�5l�V�|�j��)��?��v���        =VP��1�?��B�Q��?:q}�s��o��E�&����м ��$_�-C?V�qm~Uv=��x�cܙ=q��u�3,?�l�G(Io@^-l{�x@o����R@��ض�=�;���?�����8@>��|��?�      @/��[W>�                                A�e��@  BL+��  BL��                           >��m:Űi@��[� �n>����;�WA�o�7��>�^5%�
[A�D^� �                                                =�%�)�@w��q��?�م�����Eޱom>ad���?>��%�=�F�'���?����[X_�Q .+�L='H�5�Z> jj���>��,E�Ͻ��	���?�ַ����5 �4�S>�T����>Qڪd��^�⠄%                                                                                                                                                ;�Sט�#>3����Τ>b�
衻ꇑ�jL<}��b�m=Y�.e�r{<�V�t�*>L��Uc����
�;�?�ꢚ�<uR��i�=s�ro��<�)
��Sj��JA>����<�|���Wt�ǫ�#v>b$(�5`                                                                                                                                                �>%.>����J����8���ŹG���9y����>�I�]̳�>$����>ɝ��d�>gQ��y�>�W�5�H��<���	�����]��U�\~f�J>$������Ё�X����s�"����h�9�>�V��L?�U�W�ھ�>$��^�Zv> ��T��>:O0>���U����>5�Xp�@&\0  >-}w� �sYb��Y����vV�I�C��4�/��Ѐ&��%<@!���H  >2:eo}� ?^�s�Z�
?�H=�c��C��։L��{�"�wT�                                                                                                                                                                                                                                                                                                �Y�$� >=�>�k  �sz�Z�(�����~%���.EU��ΝD��K�Z�kt�� >@���� ?^�@���?�H?,G�6�C�"`����{�"Vx��@m�)�)þGy�{�E�>s��$�@�sr�Wm>�F8Sܣ�>ɢ�W�`�@n5<b ��L�1L��n��g�o� HEo���AS�#2�a�?� �'�fؾ A�I��|>/ΕR�
e��_�&�-˾5rS��ľ��$~Ǽ�\��8R��_��N>34�L�T�'*)�霗?�H?�ئ$��x&�x߿|1��᧡�~�[ޥ��=l6��b_b�Ih�U�(@?p����ؾ��Q"�W5�Ν.IFkA�qV��G>߷�B?^�g�c�?�H=���S@i����>;���K�DBZ�k��>W=X(�Ml�              @�P�@��4DAf$@���	| f@��8�%wA��xt   @�8`uR�N@� ��x��@V|�����@p��
d��
���?t�/�@0�G�L�BYB�L� �B�h%fD���_Ú�;A��(İ,ف����}�P�Y��d�X���/�!��{�?���3�s�        =!��q��>����*�?L���>5=Z`cݡ�%�����x�������?X�H�c��L� l~=�{[���*?$�\�4?�8Ѐ��?̢.B� G@p��
p"�
�]��Q@0�G�L�?t�/�?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?���P��~]%	������pA��l����<�q:8AH�
��2                                                >���iN���2)	|����-��}Q>"���������'��?���F���a/���k&?�d���e?x�{ý>-Θ����>�Z��d�?[���"�=�}lm'v[?���ʉ+��4r8H�ؾ>�.	�-��1�g,ش� ����;�                                                                                                                                                <�k��v־NкA4,��r�H�+�<@d"F�����[�>�3[����S��/>Q$�.���=�RELW�<�\�C��7= x^�	�=��&���0��4���>��+�i@�/ߐ�P=h��C>�z;K��[                                                                                                                                                @V�4��R�>Ѣ���"s>A?f$sv�@Iiy�5�< �"ܿ��;0@�@Q48�۩�>��� ���Sr$�F��Hn�o�@R
:�*�~?'I#��\�Y�����|�R_>�sF$������M�Ϳ�[�#y�?&�=���V�F�@���S�w!>þ� 8�q?�³ODl�Vb�R+��P����@&���  >���ܐ >��X�*��ʞ��l�9�=�M��I��Ì�s���Q��� ?{��RY'?�#��G�6@�^3�'��BoG��@`)���i                                                                                                                                                                                                                                                                                                ?���$`  ���uq >�`��r���Ɋ*Q��*��Q$�K�"�����x/�� ?{�j�n?�#����@�^5J�2y�Bo��\@`M���	@�[ةB�Z��A�1�G�?["�!��@��Ւ\���Pf^a0?������IAX�]�S'��Y{36rҿ�#��q����AR�����)����?�m{�'H7����$��>�8��Vz�?��?�����}5�M��f}S����ً��~?�y?�d�?�j�f�%�@��$����}˞��?�~d����a�Zq���Rèe�>�V(�f�@q�w�(�?�G�8V�;��,�!�����?��,�?؍�YW�@�0~,���@��h�9ؿ�0�
�(A����==+Q��+cX              @�T������R7W��@���	| f@��8�%wA��xt   @�8`uR�N@�PU�@V|�����@wl}���:��?_ ��Mb@jɤ�/������  �`��A/Dl���m�uB����'��p~�U4�PC"�DC	�D1C�zɶKB�+���?���41��        =5���4X>�����?L�M.��սX��l�;��H������(���h?'3\��n�=���`2�=�.j��F�?<'�1�Ns��F�#�?�j����z@wl{����6q@jɤ�/�?_ ��Mb?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?��f-e��b��I⿿k�L�Ae& ?�s?�+<���vA2�{���J                                                >{s��@'�-�] |��%{�%g���m	S|wK����V��'?�)�E|�2�Ķ{���9?���`��?w�����=;w�В^>cK!���?3�h3���=�����2?��("B��4�1�X��>�Ia��>�pG]�>�!y\'                                                                                                                                                <�JI�Tӱ�Ib)��B9�yu����BxGm��޾.߮=��ǫ���:蛟I��>L���A��=���%���;�I�A!��<�
���D=��?�"�Ƽ"S���(��q�i�>���C1&���Bz�?�8qe�J�|>����|%                                                                                                                                                @R[m�2�>���3<!���V5>�@J��'#t�����M�� ]k�v�@"9m��P>�<-����MKPꖥ?�B�g���.���7ݾ���يZ��T��ʌ�P�e�4��>&��.���v\��_�W�ha%>�Y������T�*8�v�d�Z���2>�=���v?��GZ7�T���WqS�~G1n,U�@&OƔT  >�p��� >�m֤����Ls�ҹ޿C�*1�"�3�H:�����+��o� ?4�;�[�?�����@�,�����B�\?�qͿ�OR��aQ                                                                                                                                                                                                                                                                                                ?�[$�   >� ���  >�[�������s��=���'3r�'>�4��r�Kr��O��~� ?4�܃)��?���ʕו@�-ԵO�w�B��l�����O]wD��@�m�!��?��Y�ҿ:>���@��w��h��X<�X� ��c��2@ݝ�,R!�N�#�rв����(���� t�w�AR�Ow4ӵ?�ó��$?�:*0PI�>ż��;��������!2?���	����7ɖ��#>o��d�n��*�h���]?5L��kA�?,�\��s@�>�"3��;*��J?�l�2�}@p�n�>>>�ڑ���8��>_`�/�@`7S��5��J��Eg��<GeT����	OU���?D���!�?����p��@�����H@�W7�n��?Z����H�@sI!3o
>=ծ c�              @�J�5�m^>e��3@���	| f@��8�%wA��xt   @�8`uR�N@���^m@V|�����@i//��:=��%�J>�OB��'�?�q%�	��@sI     ��9G��  Bÿة>�@�����)�D�ֶ�H.��]p�o�M�2t'/�:1�gA�����?���N�sH        =V��s~� ?�,����B?wxq��˽�X��<���_���C��7v0X*7?V��%�^=����=rS�ื?��6�3�@]�}���@p�	���@i//��=��?B��?�q%�	��>�OB��'�?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�(]���@�1�d��*>Ҥ�'�:Agd��>�+�M��A=?zV��                                                =�O�
�T�@�Nk�f�?���g�Խ��`1��>`����9??hF�kU�=����.�?�e�,���N�P�NH=& �*��> 
Ħ~'C>�c�l��m����Q�?A?�����5 �za��>�X%[	b>RX����X��#���W                                                                                                                                                ;�_���>3R~eƩ>S�A8���8;���<|��~UB=Z�t�fOw<���͊�>K�)e�����l)�;;��X{Uێ<t�8�e�=tc����<T����R�i"���>����U�~<��q�_��R�l��>b��5q�                                                                                                                                                �<{ ړܞ>�"�<�e����������.�����YBL>�"{��>�<z����>����;�>e��k�>��F��f�:���!����W��� �Te%�F��>$��{�:��1�Ԋ���L*�����Io�'q>~D���>��Te!
r��>$�OH>֪��&>8y�(D�F�Tc�f�>g�)lYj@&\]�  >-��n  �t����,��l�%�D�\A��c�Џr-{��@!w���  >2V?�@ ?^@5W���?��d��0�B�3�#�z�z LU                                                                                                                                                                                                                                                                                                �Xxk�<  >=�g��@ �t8�����t��.~���{׾�ڔ��\�Y��p� >@�q�  ?^@bVd�M?��f��X�B�B��S�z�y��s@l��6g�G{�U�'>t�F^"i@���p���>ݕ=0�>�"�:H4:@l�L��z־L��J���n@�\�5���s��"�AR�C�?��������uS�RY>/ɓS[*��e�٬V��5�U�p�Ѿ��<�	��)��(���x�OD�>3!�U�~�&�px���?��g����󍿅Ώ��z���֬�|�ْ�M�=^쒂{��U�#��o?ss{��h��!�mc�������������>O�aQ?^@_b��S?��c�}@��b^4�>;�f$A�Bce`�=A��f�              @��q��g>�G��i�M@���	| f@��8�%wA��xt   @�8`uR�NAbD�q@V|�����@3��>M���:K?�b!F��@$�n�¿�Bcl�_@ �+BJ�&|E)g�P �ZC��w��zDx���L/-��Լ��/�D��h\ȇ�C^�=�*[?���3�m        �&\Iya{>�������?L���1���>m�&�=���E���s΁yj�?����lr>��QY���d\Ǜ�0?*0��m:�l\�����?r��V @3��@>M��C� G@$�n�¿�?�b!F��?�      @/��[W>�                                A�e��@  BL+��  BL��                           ��1ᷢAl�]��@H���c���a&�@D�/�$T�AUe�E                                                ���l`�/A@!h��u���(?�g���p_>w�����7`?��JF��g>�2�Ǭq?���W�S׿�.]B�[U�E�A^,'�>��K����?�!6�yř��K"��?��
o�v1�3JZ�F~�������?4wP{&�� �&��a                                                                                                                                                �⓳\�f�>15(x�ξ
4֪�z�������0�,��͌e�>?/­q�=֒�WZ�$(��m���{����� �{,�=3d)�*�I>&�3	<[��Cu����+��e>��}S��=N|���(��!tR�
>�W���b                                                                                                                                                �8G�P�������kGK����`Њ@9�RԿ��j�C1D��4�Kj�D�Y��J��Կ5HX��>�)3��?��͔�E�Z� ��B�t�����@,��"�V?d���P�úbC�O�@
�K�"wC!l�o?;�J�h��RkJ�$j>�1���>�9�	ӂ?�4����R5��6���Y�N���@%R���  >��qZ@ ����p����?7��SI=M�Uer�j��}�h=��0CN���B�_�:@꦳V�-o�@��x���U6}�DTi                                                                                                                                                                                                                                                                                                ?���R�  ?{�� � ��<*Q/G���r�k{�0V�w��S�V@j������&����1���M��A�Y_��@ꦨ����@����,��U6�	=m@��#�O1?����2�s�;�zL@�dZ�O_��� AM�3��fH�fA!?�X%��?뇬.3��@;���^Bj�s�o6\AQ�F����@��y"1'%@�m)�wS?48�>�>��w��T?�⚱�J��1��IV��?A��[
|���P�Y�}A��Gn��(�+@�a��h#���5���zu��S@~M���?'��`>�>��T:@�TQ�����.�W8ջb?:^��\���eM�̿�Zā~����;Y2Ǒ@喂�>|(A���fd,@%���9p@mR�.(�=z�'��4              @��:�GK>hJZ�ڬ6@���	| f@��8�%wA��xt   @�8`uR�N@��ϝ��@V|�����@/p'D`=��=/�>�;B���?�y3�c�mR�    ?���  B�:�w���@�J���C�16���O�Ǟ��/�Ό1\��c�͵&#?�����uK        =W`��{X?�q�.(I?�ڟ��ܽ�=���恼��GB���1WqN��?V���:�$=������!=r�aG,�?�U�B\7@]��y��@q�?���@/p'D%=�#VH'?�y3�c>�;B���?�      @/��[W>�                                A�e��@  BL+��  BL��                           >���.��@�}���>�m�H}�A ��v�>�>�0|��A�P���                                                =��L�@z�y�?�E���k��΅:�"w>`r�#�?@4t|��f=��<����?��U�t��KP'�y1=%GRRv=�D r�Ի? 2OU�E���(���?�-�-PS�5VM~�>\A��1j>R�F�G��	Ҏ��                                                                                                                                                ;��ڃ>��>2���f>2�@� ���Ӥ�&<{��	��=[/���<�@>J�N�c������T�;��ſ`�<tO\.=u
�8���<��Q?ɾR�ӕ��>���?Ƽ�%�K{`��l���)>c?J�H#�                                                                                                                                                �:�{��Ol>�f�z���t���g�6������C��/>��ʆ�Hz�:��+�>��W	�=>c�����>�]�AqV�9WT����h��.�S40jYH>%����X�ϱ�90ˆ����z�=���l691�s>|����,N�S4�=%;>%�	� �>L,�O I>6�yN���S2��:>���n]@&\��  >-���B� �t������(6Y�Ft��C�D�СǰZ�@!l�;�  >2w���� ?]{r#0�?�C�t
OS�A��~0�y;�;�                                                                                                                                                                                                                                                                                                �V���]  >=�?�W  �u>��������0�ľ���R�=\�� ���H�Ws�@�� >@���<@ ?]{C��+A?�C��e|��A�M��0�y;���k@jR���G��X�>u[ʚL��@��C���>�͆��A�>ʯf��+j@j��LF�L��~��m{�k�t���C�H��AQ�M�H;#?��Ch^��Q;�{h>/��R8�Ϋk� M�5��&;C�����U8zc��Vk؟����F��>3+�U�뗾&d偼��?�C���ɣ��-=����y`�7T���z���l��=a)��O��VE��/�?u�#�%/�����̾�  ƾN��:��>�L4��?]{@{e�?�C�:�%@���2q"><1��)bB7F=O�v<�Ll�               @��9XZ�U>�0����3@���	| f@��8�%wA��xt   @�8`uR�NA
k��1�@V|�����@����F�>OD�_,(�?�R����@(�hE��B"| 4�� �5\T�|fE)C���Ѐ��22l��J��g#%�!4�i%����D�y�-�CcڰE�?���3��g        �3t}r�S>x���rd?L��E������е=(f7"���oW�'#[2>�M���k�>./�U�:��M�o䰗?�|^U�i�h�̪�=?��#��!@����F�>OD���
U@(�hE��?�R����?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?�!s{M.A�8tF@R!�Ϊ7AZ�_	��#@RH2��7AY���' W                                                >�e��@�?�#6��Ŀ����(U�>Q)� 
�>��Řg$?�lh����>���c��a?�t3y��,�O���b"�A���B">����%�?��s����G+�?��o�8S��2�~����c����?>ԛ<������o0��                                                                                                                                                <� _����=�Ʋ���Ͻ���o;l<mG�T��<�k�0�q=ڨ�1�=﮽7�>��(��V�xу7��*���F=��P�R�>��ce<�<\����$,�.k�'>���I��t=c�)����obGњ�>�i�N�5                                                                                                                                                ��@���� >�E�{��e>tc(�YTw?�>���A��?5�h>�b���E��:�B��|i>Ϥ(�0e����X*�W����<]�:�A�\-�?O���~��"Y�_���?��F�@�����)A?��W�E��I��_?�J�:�R��{�Ғ>�����R>����?�P����R���9L�C��9V��@$�$�  >�ڒ�� ��\bg8����Ɠ�$��[��G�͝�X��0�i���Z[� ��3��@��`�@�z�)�`�?��I�xp�_,��^�                                                                                                                                                                                                                                                                                                ?�k#۠  ?�Y
D ��������R� {a������V�T(Q��{�^QP�����t��`e(��@�z�?�b�?����z�_,�3�{�@�QK:w�ܿ�����,?+��ҠQ@���Ժ������s.��?��/D��A&����F?��{���6@0^L��J��)c�AP���v@o��!ay7?�ل���$'���:�>ɢ�s��?�q�����,.�?M0¼�Q��A������/�Ex!���w@��4�[����� ���Ь/3�@p%1���?
Zہ�<�>���s�@��g�/ڑ�$p��樿T����"�xzP߿�GY��O�Ri�2q�@�6E8'�@A����^@6o���l�@j� ��={Q�Cs              @��J�1xq>j��Y�(@���	| f@��8�%wA��xt   @�8`uR�N@����I�@V|�����@���oN=�����)?>�)$J�*�?��ru��@j�     ��jE`  B�9*�ҋ�@�`�^���A�v��4��x��D�+��ݱ��a7�N1�?��įτ        =W��#�Aa?���J���?}ZK��V��"8���ϼ�mF&�<;�:$A��?V|/��=��6z=s�l�<�?��x��)y@]8�̿�@r��qήG@�����=����'~?��ru��>�)$J�*�?�      @/��[W>�                                A�e��@  BL+��  BL��                           >���h9?@��3� �>�;�j6�A ��5j5�>�+�=X�AI�.�c                                                =��;�U��@O�C�K>?��&��F��6��95>_�[
�,?@��/\�=������<?�*��"6��H*)��p=#�G����=�Ӱ��? ���<����W���?�\�r2c*�5!�:}~>	�ݪS�=>S�gasDؿ��)�z                                                                                                                                                ;�J�4��>2�� �>-]?�5��%�c|�<{"��B�a=\X���v�<�_W�>J2�Z����d�i�e�;�{J�G�<sϯ�!�=u�'wB��<ّ�}���QyC���>��&��H��7���l����HK>c׬>h�                                                                                                                                                �9X3ȝ>u���eN���^�����jQ���H��1�j>�ʒb e��9�k>uK����>bI�o%>������7����1��H�99��Ro�1��>%Mٳ��U����Z��d����پ���K�� >{�H�Rkܣ`>%M�z��>
�m�=>4�TV���R\C�=)>ᤳ�2@&\ �  >-�j=(� �uҎ,�UJ��?B`[�E�H �����д�� @!a�s�  >2����  ?\�]�7?ޢ�ʴ�u�@�U\�?&�w�S_�2�                                                                                                                                                                                                                                                                                                �UX���  >=���@ �u��M���F_`k�X��>�=��c��j�U��� >@ϑ]�� ?\½b��5?ޢ���@���g���w�R�s��@hǊ�C���G�1��>>v3Nܣ��@�UJ	�>�5yٗ�N>�3PO�\@if�鹣ܾL�`a[޿l��~�=�������AP���5ڬ?���8ݾj�`3 >/��Q����3��675�LI���>F*���T�%����mL����>38MN�3�&钑w[?ޢ��z狿񬎉g���x����x�W���^=p����=S�]3d��?x���.���ח	���c�<�I���0��>l����X?\º&��?ޢ�=�^�@�I}A	><��w�B�Z=�Ǭ=��g��&              @�Q�J���r⑧i@���	| f@��8�%wA��xt   @�8`uR�NA���_~@V|�����@"�����SU����?�Ӝ��dP@0!A�GQ�T��A>�Ӳ)E5�X�b
��ȹ.��j��e���HDA�Y��D�S��@(�b�{^K��?���3�Ԍ        =5��n`�.>l8LIaH?L�@hy_!=u������16u|p�2�fUnS4>�k4�BJ�z2�؇<=�C-h�?��A�y�a�#d�+?��_��s@"����SU�$��@0!A�G?�Ӝ��dP?�      @/��[W>�                                A�e��@  BL+��  BL��                           ���O���8	�����S�[��$Adѿ�̘I�S�s��+A_�4o��                                                �J���(ɿևϔ�����R��s޾��s(੾��]2�º?�X(��1���,��wN?�w�P���rͷ!���>,e���4>��clW�?�p�q�>=�c��̧�?�^�!���1	P;�F>�A:Ԉ�]�:�|=��1��͆                                                                                                                                                �f���,��xϾmȽ��wQ�C�,jJ�(C��E�j�PE=���&gսg���U<> �"�b�Ľ�m��I��<�r9���=��U��h>�d1�g�`��w~�����R�>��%E�+�qf��O9=��3c��>�@r�"�                                                                                                                                                ?���^�h�/l����8�@�Jh�?ʙ�Oh���Ծ�Z�'��&�"������)�����r�b����/��q�&db;+m>�vj3Z��&:�����"z/��U>����K[�?�l@�����i�=�?���L�b�R]��߿�uos��w�T=s?�����{��RVRk�y,�=y���O@#�y�<  >���Ԛ� >�=�؜������y�e�����]��6/��� w T�?�C�HR/@.�׀78@�'�~���<�i�f@Z��Z6�                                                                                                                                                                                                                                                                                                ?�[*�  ����Q� >���+��������1�� W�?���\��r�H� �h>?�����K@.ϖ��j@�'�*��<����@Z�}��O@�3UZ9�࿅�����n?��#@@��bd��s%��i?��[J�A0��T4�'�/�X�~���no�+9ƻ�%�NRAOW��,���m�MZ�?�w������r���@>���Zg`�?d��8� ��f95k?3i�Y��ٔ���@,�����@\�����@�$�s�)�b�^@�{n9%@c�n�2iI?\�ydBz��b�?(@�<��~���</RyܿX��NԽ.�(��BL?��rĽȆ@N�L���@�1�?]��A ���>���?O�Nƣ�@{)�A��=�r����              @�T��i>m��-��@���	| f@��8�%wA��xt   @�8`uR�N@������@V|�����@$lkmb=��
�7
>����X&?�H6LΦ&�{)�    ��%t   B�����th@�A�\(��@~ g2�F�����lN�(	'��D�]�Y�`�_?���dg�`        =XoW�<?��m(*?����ｯ#���˼�
$q�s��P����A?Vi�8�Ot=���!�Fe=t/��E��?��*	��t@\�=��LU@s����
@$lk,#=���d�Uf?�H6LΦ&>����X&?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�c@kw�@�<F�hd�>�G�AFA (�ϙ�>�TfeJp�A{=��jf                                                =�'�,�L@��L[�s?��\(a�ֽ���u�x>_#q���?A4��p��=��.Q.�?Ӛ�I�
m�EMnك��="�d?Y��=����~�?2�7��G���Uրj?٘V�]7M�50K�~�>��쇲>T!d��?���:�\�                                                                                                                                                ;��?�i>1�mLx�>}�
-%ػ�d�ߖr<zj�e"�=]1��z�<�B�Uka>Ix��x佻��E�ǲ;���mB�<sXJwS�L=vWo��	�<lay�D�P����.>��9�ϝӼ�Q��9�V�ʯ�V��>doˌ��	                                                                                                                                                �7��O��E>b���������}@��z�ݾ�)_��>��Y���7�M���>b&��j>`���4�>����ĉ�6Z��g��1��?=X�Qdf�ڶ>%}i��t��l��""��������]P^�>y��a�!�Q`��>%}_0rW�>� 0�>3St/���Qmù �>�$t��@&\�J  >-��M�  �v�e�
��������(�I����M�������=@!V	�  >2� ��  ?\��?�'���I�?P>�@��v�u��S                                                                                                                                                                                                                                                                                                �S�
�� >>U,#� �v���0�I���e�V]���ݣ5忾ϥ�o�1�T���	� >@���  ?\�Ǐ�9?�)�B\��?P�j����v�u;�ެ@g_���G��6�2>w��S� @��[��>�����>˯�u��V@h fe`Ҟ�M��qGq�l=C��6����AOP�� ?����L�]����L�>/Ѣw� ����k�v�6�VE�r���ݨ�[:�u�C_>n꾜��Q1>3GH�UL(�%�NQFQw?�*��\��ڙ��9Ϳv�lܟ˿wf����=p.�=>Z�F��T?zblq]�F���K>�m�ϥ~{�gt���&�>�O:`?\�i$З?�%��>@�	��L><�ԕ2��B������=9ja	rS              @��5��|_��P6@���	| f@��8�%wA��xt   @�8`uR�NA֩{w�e@V|�����@��d#뿾���{#D�?�|Qs�-@5�7�&B��*��BM����f@EH�u䍳L�̑��
pt+�sDw��N�D��o&��Î�Jg^�?���3��        =[PdQ�0=>Z�Կ���?L�W�ǎ�=��h��''�\e^HD��[������>�Z6 9� �5��o�=�����%>�>��+^�T\�-*cG?�l�7�
@��d#������q�+�@5�7�&?�|Qs�-?�      @/��[W>�                                A�e��@  BL+��  BL��                           ����9���<A�@�!�����2��Aiρ��{���
I�Ac���2}I                                                �oB8�ʿ��2-�׿�L����5L Ȑ.W����&�?�,|���:�JQ3�?��
��ʿe��I*>3�ߘ��
������p?�����>i>8�`�a�?���S�e��,�AI�;9?-FDW�ڿde�o ����*�                                                                                                                                                ����d�h���Xk������̓� �R��@����6�v;=�ϠjzTk�7������>(�� ���R`#��(<���j�vX�r�l�1> ����(v���ʶ����֤ϡ�>�(�T����g[2!�8=ڊأ�>��� ��                                                                                                                                                ?�Y�@�����N�} �Y`�vn�?�ޒ^��ʿ��_��2���Q�֦��A���fh��a�?�H��3+��w[�H2��C?�+�|���k�>��$_Hr�<�?+~_̧>���Q�K�?��Bu���%�\���#� ���M�R1����8�6_I����&�$�6?�=8�(49�R�x_�!�\K�ks2�@"7Ȉ�  >��^E  ?��"�Z����O�e�q��W�6��a��>���'m�e7p@'������@Lk@�t(�A���hN�:b�ݗ�@��;��V
                                                                                                                                                                                                                                                                                                ?��   �>��Ke ?3b�?����ѡ�5�%�3�/��b��x�'nt�5{r@'�f2�2@Lk@�#�(A���۪�:���@��8���@�z�4]h��>����H��E(�ư@�/�uPʿ@�_.e�<�⡇:�]�A8�;YFp�j}���ϡ��I��/B�%��%�A�AN���
1�Â~�<�]���9����?@��X��}��& �ޖ�p�tś$�'��~d��?q�[(c��`8��҅@g�mUf��@�H���(lA	{k��M�!��7�@���ܝl@Xp���?JW·ɜʿmEa�@��n�U��@�}�N��U�W��'�+����<@,	Je�)@$��u��S@�&Df�i�A)��R��{�sB�Ӄ~�@Uāj��<=j�Ӊ�P              @�)kx>p3.jL@���	| f@��8�%wA��xt   @�8`uR�N@���M�. @V|�����@�q��=��J��ѫ>�*]fT?���C�܈@UĀ    ��l�sp  B��U�X�@���جB�>̈́�����V3)����%^��t�Y�N̊�?�����l        =X�J�{Z1?�|��ԑ?���lֽ��^\q��|	LwX��s��H?VU�@b��=��}G�m�=t�l4v��?�������@\�>]���@t�w:#@�q���=�������?���C�܈>�*]fT?�      @/��[W>�                                A�e��@  BL+��  BL��                           >���s�,0@�U����>���"��@���=̻�>�I��b>A�+.)                                                =�w��!�@
*G?���$�PY�Ͷ,-6},>^Ym��Z3?A�:>���=��YԿ?���|��B�}�6 y=!<�)g� =���I��?�?�,�~����`T;?��Xu��U�5=��FM>^vb�*4>T��؜��B��
*                                                                                                                                                ;�Uߏ(>1 c�5��>�
!��2��5(Qh^"<y��^w��=^
a;.�<:ī"_>HǸjC!���H� ��s;�d�u�m�<r�XA�I=v�`N!�C<]'�,!��P|h�[4�>��K����wd�����4:��>e��@L�                                                                                                                                                �6PC��|>S��צ����)`;.�C���qݾ�$��G�>��'XYf�6O���->S���>^�!^֔�>��(#_��5)/`2*׽�8!X�P4pU�R�>%�2�~����|"�N0��n� Y:5��`�EoF�>x| ,Ŏ"�P4l�*��>%�(�v�><N#�sh>1������P3��Ck>����@&\�"  >.!�ͅ� �w�	jԠ���4Mb-�^�KWy�^C4����!�T�@!J�  >2�u�n@ ?[s��&
?݂�����=�bL�w*�uht�|Ft                                                                                                                                                                                                                                                                                                �R�� >><�Jx  �w��:�\���:I��ľ���~�t���I��A�S_��  >A'w�` ?[s��g?݂�BD/:�=��Ddj�uht)L�^@f�m&Z�G�n���^>w���\@�F$��>�|@괄>>�%��$�f@f�'�.�ԾM,
���ks�
oP0�����*s�AM����?�!��:o�6��-[l>/���eJg�����W6�7�-��L����y�����$Ƙ����x_�B9Y>3X� ����%c2��T?݂�B����M�wr(�u�3���vE0���=`D�D8�J��^=q�?|��AS̾���_8[���8�����JJL��>�	���?[sΎ�t�?݂�ylu@D���#�>=K<{m1B�+����P<���]��              @��!�dS���𾫘&U@���	| f@��8�%wA��xt   @�8`uR�NA �.;0Xj@V|�����@B��.��5��ψ�?��ɥ3�@Abщ���uP2�}'(KV�g�Eo}֝7�6�<˴���D�����mE5ᷱl�D������#<e�gj?���3��T        =�g�rl��>9�����a?L�g>��!>��
Wǐ��C֕��P�D�\�I4�>�Aմɿ$�������>���`7��>�uD����;��[�?��)�/�)@B��.��5�����@Abщ��?��ɥ3�?�      @/��[W>�                                A�e��@  BL+��  BL��                           �tZ]�	��5q�,GZ���p�x+Am�Vx�޶����X��Ag!����4                                                �fwr��é�⭿N���J=��B�5x��>�l��n�8?���u�U�G��N��?��8�a���S��{;�&��g����?����J?�3�|�>�>�P���S?�[[�[���!;���r5?�z��%�ӿ���D����+�40                                                                                                                                                �$����Y~�஛��	h�jH��*c��w[i)u<�߶8M�3=��������ZF�>&�����~n�a��8槭n�> �WZy�{>2Q�{�c޽9R�8������#V>��6��6F�7+�h�=�>a �Dk�p>��>���                                                                                                                                                ?�EF�@K �$/���ܠ��6t�yVY?p�ݾ-������k�1>ٖ?��V�ۉ����@�r��uhc7���I�0�xf��q;��V��� �sA�
�F�o�u0h���6�4F�@(,�pV�?�?h���7E83쭘@?!X��@�R�]:���Ҙ�/��i������࿳%*�J��X��M��X@)�ȮF�@�@�  >½��   ?��m q������h�Mӿz���l�e?�����0�q�� @����@��N4�fMA�R�y�7�����A?���                                                                                                                                                                                                                                                                                                ?�xkm�  ���g� ?��	`ĉ���xCB}��7U~�B��@9�;��>�0뼯)��@��:�g�@��M�A˸����7�"@{��A?l��~@�|wSƾ���51�r�����y˨@�Ϝ�+�@�1w������Ỽ�UiAC��̷9��	�\�@���$cg�S+��6�K��APU���>f"�4Bb�)�[e+@{*��� ?���a��_?��v��B��� �@;���i>��~>?A*ۼ��[AS#a:>]A���¹�1�v&R�oA7�n�Fy�@F)�r:��?�mZ3�w���)��@�W�T�@Abv�#���v��� ��$d
@�4W4�+���Em�Ê�M����A6�6�4�
�L�1��@�b���=�66@              @���Zl�8>q����@���	| f@��8�%wA��xt   @�8`uR�N@��J���<@V|�����@阉=��@���>�&44�?�Y��:���b�    ��c>*0  B�Aa@�H�I�ܼ�<ؒ���A�� 6��9�"x/��K�V����{O?��FR�        =Yp�
��?��9˒�?W/�����`��m¼�9G�
Q���p�6�?VA7��.=����O�=u_S�&?���U%�8@\"�8�Q@u�%h_�n@�%;=����r��?�Y��:�>�&44�?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�O�ɝ��@�&WG��>ֽ�|�@��(b��>�AW�f�A}8&�G�                                                =������@vx���?��6�q��̓i��>]��v��?B3���=�ng'�v�?Ғ��ÿ@O���= �c���=�y�C�!�?1��1�����X���?�0�0Hx�5J%>(r�?t>U]��O�{��O^��y�                                                                                                                                                ;��ۿ9b>0�.�D�C>?r�����
���<y b���C=^⃛���<р�̂>H!9a9#���/�;�y�u�<rQ��r/=w���<<���Ϙ�P͗���>��[�D"���������R��׿�>e�d��Z                                                                                                                                                �5��C>I����O��d���=`@d��8ޘ$0U>�kd�=�5y2 ˦>H��G��>\R��ק�>�Ǜ�I��4n~L8`����J]*0�N����>%�D�k����J�O4����,���ۍ��?���b�>wSX
W���N���՟>%�:�S֦>��>A�>0���r@0�N�<�V��>�����@&\X<  >.FAM�  �xv붼�������n 4�Mk�.�����s1[
�@!=�I  >3F�<� ?Z۲m�&?�d���F�<r�	�t`�H�N                                                                                                                                                                                                                                                                                                �Q�?�@ >>d��u  �x��15i����rI�����=���
x��R;�4�� >A&D<@ ?Z��
v�?�f2��h�<j��t�t`��>�d@d��o�;��G��Z�&>x�/�H@���x�>�Q_�_K�>̕���@e��6�`>�MW�Io��j��+J1��sݯ��ALlq1�?���� [о�Zz @>/��)��8���j��7�!��v?����$��p�`�0�N��2܌>3k���%X�l��?�g1)¾���҃r4i�t�=��UԿtȭf�n=f�S�hܽ?��:�0?~���'E����-��C���4MP�{�?�3�>Bȣ}�?Z��a���?�b<�� @v�䅔;>=�E�|��@t���)�=�K����              @�ZΧ�'�>sZD��+�@���	| f@��8�%wA��xt   @�8`uR�N@��]�yƅ@V|�����@�A7W�=�D��
��>��x�0�^?��r��e��t��    ?��   B�ȱ�80<@�p���-��;.�"�����Uj?�� J���?�S�+�N�?��q�*M        =Y�!�j�F?����Kq�? ��4[br�������Ӗ�"�p����㣾*�?V+�IL�=�Ƽ����=u�{B+�?�я� �@[���:"@wx����@�A7W��=�Dە5i?��r��e�>��x�0�^?�      @/��[W>�                                A�e��@  BL+��  BL��                           >��_"�v@�ud`P$>ם-r{�D@�C���+>��u���^A	��'-�                                                =�&S�C�@��3��k?�q���]��]=r��S>\�$��v?B��_��=�Y�^���?��W��<?���5=,�kl��=��:Ѧ�?��2����0����?׌E��/��5UG(Lr>���G|�>U�\o��f���I��                                                                                                                                                < ?/� è>0�qR�`>	� x�Gڻ�����<x���^$�=_����<j@��RV>G��8����Yn7�Q�;���dJ>f<r����=xG�¡�<Ʌ$�q�O7S�d�>��j��m#����0kn��)*�*?>f6[�V�                                                                                                                                                �3��콋>B;}:l���j�{<�8Ă#��b@ݺ�M>~{�6r+��3�b�X�>A�C��&>ZE|j��>� 0��(8�3�)����-�6@�M.��@x>&gR�ꇽ�ƹz�T��%�M�1��5���>vBS;���M.�핹 >&\��T>.��JM>/KM~����M-Pײ> ��~e@&\Đ  >.l�9� �y]D����F>:&z�N��=�����U��U@!0�n�  >33�n�� ?ZM+;}^?܋�mĪ�:��Q7t�sm��E�                                                                                                                                                                                                                                                                                                �P��!�@ >>��~�  �ywQ���f��KU�=��LM����2���>��Q0��� >AE��;� ?ZM'���W?܋���;��:�5���6�sm����~@c�cņa��G�yES>y�a$a�@�U�i��>�Bg�u�c>�W���@dz�#�)t�M����>ɿjMH��#�����oHAJ�70$l?�K�<	uF��=��5">/�jSڙ~���$z�%,�8\!	���Jn�<���A4\���JRR%�>3�LH64�$܇��5?܋��������@7�s�:+����s�gk��=^�[�-��H��h�?�Z�je`�����n��2��U7����Y���>�2�#ܰ?ZM#�6��?܋���o�@����l>>��г@NGH~
�=h"Q�x�              @�ǔ] >u�z]�@���	| f@��8�%wA��xt   @�8`uR�N@�����@V|�����@	�w��=ݱ��ҡ�? y���*?�o&s�v@NG     ��\{�@  B��z�\��@��F����9�Z��g���1����"z���QzF�Y��?��$e�=        =Z$�J?����6�?!c �K���Je�U�����о�G���M?V��q��=��(���=vm��O"x?��~��#@[]��qخ@x0=Ĉv@	�w��{=ݰ��H�k?�o&s�v? y���*?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�Q�a�@�4��ӌ>؀�z��<@���U��>�S�E���A��;��                                                =゘�/�@i�t���?��Ys�߽�>_��U>\Kr]/�~?C1?���3=�D�׻��?ѧ�CI�8<�v���=�k�'��=�S�O=b!?/e;&;��� F�?�𡤤(T�5_���>u9\_�>V���;)���2�6k}�                                                                                                                                                < �wގ��>/>Z����>����^N��τ�=��<xj��^�=`Hs�l��<$�t�M>F����̽�|���*;��ݶ�1�<q�)�GB�=x��=u<��PHľNi=��>��x]�t{��$��q�J���lj�'>f̘2sV                                                                                                                                                �2���ߺ>>_%A�J��C$��(��<���t�����#6.>}�l�q�2��ѯ�>=�ؽ��>XnpfطW>��>���b�2P�6iJ=�^�k�60�K�KE���>&=�R�P���H�J(e��Sx�S��A�x=Y�>uF��Z�3�K�D�8�8>&=��v3>�P?�>-Q!����K�d�(> {a���@&\2�  >.�퇢  �zD���"����,*��Poy1̹��S��&$@!#��0  >3]`�$� ?Y��!U�?�0h��9b�;.�m�r����I�                                                                                                                                                                                                                                                                                                �O%=��� >>�춃  �z^]]v����v���}��Ȥ;�4���Q��s�P9��b  >Ae�@Ǡ ?Y�7,���?� R.{��9cڈDѿr��a�f
@b��[=���G�Ǩ�P>z��&ve?@��3�ٴ�>�L"��.|>�h���2@c}�X�O�M��~/�7�i�SA�lԿ�.��~AIcLK=-?��r�xpR���6�e�>0b�����e>�}���8����ĸ��Ȥ8��뼓u;I��2��8d0�$*>3��;��J�$�3�'?�!M�/
��e�>g1�r� yd�r��� ҽ3��g!dl�c�=dPp?�Y������ʓ=�f���Q�"%eG�㮕h\> N�fR�?Y�34�K?��A��@��B�D�>>��W��B=���I��=���5�              @��wW��d��᫺�@���	| f@��8�%wA��xt   @�8`uR�NA];׳�@V|�����@wdh\?F�h�0���?�"�ϙɾ@#-@���pB;VP5�] B&�`(�2_E�G"�ND)=5n�[D�uj�D�Ӌ

PD���6��HC/���?���3��        =F�`�T�>��:�E?L����Z��*rü��'�Q��urM�k? ����=裧N�e=�e�y�?����f8�i�\K�(��'��$�@wdh\?n�h�/����@#-@���p?�"�ϙɾ?�      @/��[W>�                                A�e��@  BL+��  BL��                           ���S���e���@C�)FApo$X��z@B���ܜAUCy�?�W                                                ��C�'KJ����sB�?q��BW�оl�Lځo���歘�?Θ^`��A>o��b��?�8�0 E�}˗�\1Ӿ)�u?�]̾�EW��xa?������>X�I���?�[|����3s�v���>�C����?(}�/����Tfc�                                                                                                                                                ��1+�Qo�0P,b��=��gQZ.���DQ2S�Ӽ�ow�lY=�����{<�Ľؓ�>8��eL7��Z��uΐ����5�cm�Ch�-��>E:m]���v���!ٙ�"!��	Z�>��
K=W<�'�k�O�սw���u%>��Ba3B�                                                                                                                                                @2��ѱ^��|_��$뾌�4������4G+0��C�v�����!p?�`@3R&y�����4е�Z�>iy "�� ����q�`�@3���l+>���΄��=��a��>���w\��B�n��?�硕a�;���gm*O�F���ôV�LK3{g>�R��:|�T�5��?ȁ#:2��L
!���?W��޲Tg@%tq�
  >��9�  ?=4���G��S��K�7�P�]8�P�]�bd���Ǳ[�?x���,�?ϴ�Jj=@گҭ�n��7jC�Z���'m���                                                                                                                                                                                                                                                                                                ?���@  >�1C"8 ?�x��2���P�k�y"�qg�D��\qB:@�����(?x{*b�9�?ϳ�&Kx@گ��]��7jgw|QH�%�Yܥ@�X!�gB�?轜]��tl�jp@��}�r���\��r�Y����7�t�A�.����?�v���@	��S?j��̇�5�AG����@]��@ݬG@[�_(P?[��v/�t�h��?�a��n��_L/V��f?�Ӎ�K�����f࿯�[��lR�����%�@۱�@ڒ��L}���7�Y��Tr=	@n`TxTl�?0X�"]��U���2P@�SY��`(�8Ks��v�LP��[��P8b?��xhӺ�?�rn�3f�@�Ft5E��AD~N��P?����`A�8�0�(=Ai� �>�              @������p��D�K6�@���	| f@��8�%wA��xt   @�8`uR�N@�K�i�D�@V|�����@wv\%0�&nu�Q8?pH�O@�z� �ZA�8�g�@ ���T�D~��պ%RB��:[��HĄH�����CX>�n���C�� �l�P���S?���3�%�        =$�
xX)>�'ٸ?L������= �s�Ž �SW��6Y~EA�? 9����23'H�=���m�=i?+O�p��F���?�?�e�X�@wv\%2��&q���n@�z� �Z?pH�O?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?�k�97��h��&!U���%�3~AnN2�S�J���Qw��AD�e gT                                                >c�h�S�'�r	������6H��3��/����"��y�?ȡ�<1�;�`}�}�?����}��?q�ٿ��=��,Y ؉>k���x�?0ީ�yd=���_P��?�A���3�4��|�>�Z>��o���׆����m�R�<w                                                                                                                                                <�%�~��ҾC�j���"K�	����P-�M����HkH��=���<Ŷ��y��Kn>H�=��\Z=�6H�?~<�'��6<����J�4=��	I�5+��s�z�"���u��>�`���"!;����=!$�U>�.;��M�                                                                                                                                                @G�C7�n�>�I�Q���`)�oK@%������2+4\��2�r�a�@@�A#�>s�F��ꢾߛLO-[I?���9�N@�Y}�vX��=d�cA�M�?�ྒྷ~�@��>gg�j�Կ�H�z��տhy��ȵ[>�@�Ū%�KS\�2����4 �>�=��)N�?��/��G�KQ��'�����;�ސ@&'�f  >��V�� >�S!Ǻ�`��-=<�i6�.���&�ƿ@/��+����s����?X%'F֮?�8ޘg�@��s>6@�8a�?�ıJ�o                                                                                                                                                                                                                                                                                                ?�/�XP  >������ >��Y����#<=�����g"��@��;G���w�&�?X$G���?�����@����ko��8���J~?�ĩn�bX@�=����>��*_��&����@@�g/�ˬ��J}m��O�}�@������r�Z'�¿ڿ��q���ͱ�ȸAH0�5���
��Bp@?��	I��4>��e,0��硫Z�S?~���ؿ��h�P/>Z?�ފ�~�Y� #��F?[�ږ��N?������@��t'W���ʛ�es�@c�х�﷢�&r>�X�㶠�>�@�1�4�@^�X���R��|sM���@ъ+Q4 ��]�2֓�?g��3�?�#sI�@��	��@���h�@���g-�w@g�@E�c�=��i�              @����>v�:"n�@���	| f@��8�%wA��xt   @�8`uR�N@�'h���@V|�����@���>�=� �^��}? ��B�?��.r�@g�@    ?�����  B�mi���@�� o���8�vd	W���<��X��X����N�yP�D?��3'^�        =Z��L�?����L��?"E�dDw��qS^R��Ԉ�c����k�Ჰ�?U��b6�j=���[o`�=v���V�x?�5����@Z����VH@yPe!���@���p�=� �3��?��.r�? ��B�?�      @/��[W>�                                A�e��@  BL+��  BL��                           >��s
q@��%��[>�j�B�;�@�>רl)>����nt�A83UI�d                                                =��Q��~@����
?�~�K;{��'�qT�>[��|�N?C�l#� =�5��|�?�:eL҇��4��-� �=#��Yz=�����M?��������1%�=y?�]X!'m�5i��G>q`��18>WJI�"�L������%                                                                                                                                                < ߇�"q>.nK�]5>S�����L_��<w��S0=`��=�]<�~.�>Fa��f+���5���;�U �C�<qi2�k�=y�]B�<�r}���M��=2P�>�؄�ܻ��rڬ�������>gb�F[_�                                                                                                                                                �2��a�>=�������ˋ�����,�߾��7t�}�>{Ă��O�2څv��>=\^0bL>V�ևUe3>�Q#G��1BӵR�=�h5�_���Jo�O�s+>&m����Ӵ�?�x���v(�ƾ�`���>t^E\���Jo�?�U>&m�Ny��>�͸���>+���)���Jndw�> �z��PZ@&\�`  >.��:� �{.e�A�@��q*U���Qn���R��1��0��@!�~  >3���@ ?YIS}��X?۹��� �8-��a�q�8�
�                                                                                                                                                                                                                                                                                                �M[��  >>��a� �{Gf�g����ud���ؾ���V�0���q-��2��N�vpy  >A���q� ?YIkO�+6?۹�FA�8.&0` ��q�8P�&�@a�e6
��G�
�8Ҵ>{�C�e~@�~g�J�6>�k��D".>��r��:@b��g��M�߀<3 �iI�	��a������8AH.'��-�?��љ�2��h�1��>0J������|z}m��9@[1{����K{�:<��Ps͂��۶��D�>3�O� Ծ$o���?۹��;���S*ެ;'�r"���)�q̳[Ǎ[=Y�]�2�w�R�b�`�?�T^w��.���Ɍ�/m��q&����_�:��> �G���?YIg/��2?۹ p�=�@�aT\4>>�\����Aj2�F���<�%�z ��              @�K��H꾬����O@���	| f@��8�%wA��xt   @�8`uR�N@ڻ��`u�@V|�����@��rΨ�(����?[SC{?�;�)&�q�h�:y�  �O���DUjD]e��7~���\���?&H��^��痋qD�Bك�Bc����0�?���4dP�        =8��.���>�ŷ�x��?L��:����a�Ov؇��^�&F������?%5���F=�;.��=��VA�J0?@>靜vT�����A�?�$�`��@��rΨھ(���=f?�;�)&�q?[SC{?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?��C��t��Q���z�[�Z�[+AV��g�Z:?��C���~A1�Y��R                                                >w���$�6$Bz5�#��S���o�cz�̒��Rl�7o7?Ӈ̃^�������?��pq?k�캋�/=q��m��>T�֯+P�?.}ʽ�=�~>�M`?�3�އH]�4�+Q�>�V��"�<>��;^겼��D���                                                                                                                                                <��3t>ӾAp��O�@�9`������╶v��{��s=��其�6��8>F6[,$=�&[�;�Qd}ɏ�<ʬ����=��]Yɨ�#�u�"�Ⱦ#[r�F�>��{�s����,Lqr��4�����>��V�|�                                                                                                                                                @D'{����>��.�j����M� ]Z@CK��3dH����]¾�ԯnb�@)RD�~�>>���zl(��V���G?�O��l��+.?��'>�L�65(��I�Q�X�s�V��E/=��x�/Կ��`%Y���:��۱�>�ҫ��]��IorF���Vf�v�"m>i0`�'�>�h�L��i�InXC	U�k�aF;'�@&R�U�  >��L*0� >�<k�o_��	�bA������f�*��nY�@����W@ ?��	7`?�0+��@�n�g� *�7�H��#��B_��                                                                                                                                                                                                                                                                                                ?����  >�@�e
� >���)���������m�햪�+�޷z{�����y� ?�q�� (?�/V�.@�q�[���7 ��l���B�y�@Ҍ{j�j�cG���W�?Z�  1�t@�Ͽ�$ ��K�O�|?r}�|/@�-X���V�Xo-�`ڲ��]�~ܱ����V���AG&�}<pJ?ܻ=�?�.��b"��-�&���>�ځ"˭?��H��j_���A�8?P�;@;�ߝl��r?������([��@�w�e��(���, �ɿ�o���6`@r�&���>�
�B����IAa	@jn�/Y��#]����3�������;��z��?*~�VQz�?���6E�@�d�Vmn@��& ��?K7!�w�b@i��N�1.=��Z��Z              @�Z9x��>xϋ�rR@���	| f@��8�%wA��xt   @�8`uR�N@�>h*�&!@V|�����@���M��=�z��^!�?vR*�l?���L7sv�i��    ?�պQ�  B���}�@�����j�6�mTo����
%����� R0�KXu��%�?��@��z�        =["f�7�?��1��1?#-^��4���Q���'��6v�����~i�?U�䀜= =�ݎdG�N=w����H�?�v�s�\�@Z�T㳸@zs$U�:@���M{�=�{�i)?���L7sv?vR*�l?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�g;�n�W@�by`�>�XQ��7@��RSa@�>�����A��mըK                                                =�F���@{~d��?�0��6������wŤ>[$y�')?D-vyW�=�& ��T?��\T�G��1$�D��=8i
�ì=�P��_?+P))��������?�����"�5qŚ#s>t�+A�>W�_��~����gS                                                                                                                                                <3����F>-��a�
>8�];|������X<w-�L��=a ��6<;���!->E���V�Խ�Eo�J�;���QP"�<q{�5��=z3�s�<7��C���L��лנ>�ؐw�G5����Wv����""�Q>g��|�m�                                                                                                                                                �1'e��>?�~l�d�������{^��9����)JV>z�����?�1&۹8��>?N�vy�>UH蝫��>���b��0v�8���=�1�>���I6�;��">&�W��Q��c��lg���2�#p�ھ��
�X�>s�h{G&q�I6�3}v>&�MN��>Iy�XД>)�F&q/�I5�;��f>!O��_Y�@&\�  >.�#�� �|
�	���b��l�Rw�[��M��H��ÀP@!��4  >3�� n  ?X�'u%�w?�[���	�7��0@�p��u�?�                                                                                                                                                                                                                                                                                                �K�i�� >?�7� �|1|�Q�r���c�N��D�caK�Аa��|I�MU��  >A�$�� ?X�=�ZX�?�[��*i��71���M�p���K��@a�&��p�HNOU��>|hݦ�]�@��h�N>ҟ#	Q,>�-1^�^@a������N)�p�K��h�Qq,Cv��\�.aAG3.m(?��G(PTN���0)�>0�ָF��⾚�x�9�ܵ�rھ�D�cqG�<t�Ndľ�CNc�<�>3�6��Ȟ�$B�W��?�[��U��V�'b�qP�g��p�pL�U =D��Gތ��XO���?�K�����F���АZx��&�R���m)>!>�TM?X�9mh1�?�[�>��@N�Uպ>?mF�D�BA�c�7|�<�t���O              @���q� �>��M'�O@���	| f@��8�%wA��xt   @�8`uR�NAN8�ܗL@V|�����@fvG�>Oκ�y�?�O�R"@0�i.6f�8ỪaF �8�Ȇ�!�E%��+��g��K�]׵�������DA��e�D��tr�Q�CN7�)���?���3��        �!��R�!0>m���H��?L�FZ�[��l(7�>W=|I�)�^�d��4�0�>�v����>�� �x��f��t�O?
5_Ӂ�bHB�?M?��R@�&@fvG�z>Oι�-�@0�i.6f?�O�R"?�      @/��[W>�                                A�e��@  BL+��  BL��                           ��0N͉AA>�ӳ�T@Ec� C?A_í��:@D�m*g�Aao�p�                                                ��:�ƌ��?�^	3���AnrEv�Y�z�n<)���D)I�?�rB7n�>�����3�?��Zs����p��B��%��O�>���A���?��:��R��exb#?�S~��0�̺K����K:?/��͠O����e��                                                                                                                                                ��P���=�Ž�&�/����'�u��V����G/=��X�Ov=.�Fmto>��d���屦q�k��=���="��
*X9>��k�(�<[Y<�J��!sƔ1l>��S!��=Zc��u׽���s�>�N�,�^                                                                                                                                                ��Xawp����˾�R�w���'?��,`a��?��bV�.�W���:�H�V���ف^��30>�,�U�%��;~�'��;36݅X��S3��Y���Q��x?�6{����
�_�?�~����LC绯�?%��E�u�I����:�>�ߏβ{>��Ʌ<&�?����W��Ia�=�K��LY�KĲ�@#�
�  >�!�],  ���"�����P�6۩�g�����[�Y�f�ߋ��<Ko� ��|�lm�� rub���@��(�3�������I�g��                                                                                                                                                                                                                                                                                                ?��x@  ?�(! ����)�e��N�-��7��%��X y����=}��d��{�� }� rs
�1i@�ϻ���3�/�-$Z�I���-3@���U���� L�a�?9��E�[�@������o�g�	�?�����	A(�b����9���S�G���<���u����AE�����}�g�]�?��&Ny?�&��ܫU>�Ճ%��t?��#h��c�`�Y��7?@}������K�vH_@�2 #!d@9�<Μ@y@�0%EN��lN�kj@��b�w�@bVwK�@۾Ŭe�?,>�WZّv@��6�vC�
���[�QIĝ��"@��Q��E�s6dx��=_7�V@�6Gbf�A(W���@0C�2ꃗ@q��ǤP=��;9m�              @���x�g>z��@�bV@���	| f@��8�%wA��xt   @�8`uR�N@�V�Բ@V|�����@pfqEo=��N�Bm?��0��H?�C��@q��    ��i(i0  B�2�Ѹ:@���� ��5����?���&'�!{�{��,���HNX[ M"?��Mǈ        =[\���;?��^�|�?$>��m��1u2�z�Պ^O��t��@Uni�?U�qo�9�=�� �F,=x���#T?��csa�@Z)����@{���HE[@pfqEɇ=�绹�0�?�C��?��0��H?�      @/��[W>�                                A�e��@  BL+��  BL��                           >���⦗@�f��F>�K�<a��@����p]>����AmeX^                                                =�n�uF @T���*?���ߟ��	��v:�>Z�@=���?D�;���6=����?�q����+�؏m�=���|�H=����M�?�y��K���qd.8`?�Mz����5y�uj�>�A���>X��dUݿ��׿�G                                                                                                                                                <�N�2+>,��;>3&QE�v����	}<v�!��{�=a�J8�b'<پЮN!>E\ç���/�E��z;�]ţ���<pʰ	N5=z�iG,w�<4U}�%�L=\:Xd�>�؛o���-N�����Q���}r>h��F���                                                                                                                                                �0Z�G�
>Cʩ%H��U�Q�	��M�Ⱦ�f0�7t>yv��.��0Y�Q�7>CBLd�2>S��ڎy>�
�kT���/r����=�&���(�H�����>&�[}�F�����d����7�s@����+W�>r�u�_��H��^>&�PV��>\lԟ�>(r�UN=�H��f.>!���@&\��  >/��*� �}�q�O2��b�lC�/�S��Ū.C��`�L.e@ ��P  >3�W=�� ?Xd��?�zS���6�x<�]�pN��4�                                                                                                                                                                                                                                                                                                �J*�e  >?>�R6� �}�Jw�\��j(��8Ⱦ�����C5�Я�{C���K��-� >A���	� ?Xd3��7`?�{g�i�6	Y��d�pN� �N@`KF�Xb�H*��$*�>}V-�:�@�y��1��>�������>΋[�Ƥ�@`���J{�NfP���l�hdC��hu����7�AF
�u�?���N	��yZ_Q�>0,���+ܽ��%z��<�:���3Z����ף��<���
�����q��>3�@�9�̾$LAѮ�?�|a=����l��9 C�p�L]̺ �pC���4=a����H=Gh�/8!t?�Ac�0L���>72�?�Я�6��+����gz>!tѻ�s�?Xd/K	@d?�vr�w@���l�>?�ce'�sBg�h����<��{�r              @��=v����ۑ�=��@���	| f@��8�%wA��xt   @�8`uR�NAg�E�^@V|�����@��J���b��aa5l?�x��Ҋk@5� eU�Bf�(��{��J�����E4�bj:��C�ED5t;���7���uD48?U�>�D�vM����o�w�m�?���3�y�        =D Ou�>_l7��8i?L�X�d��=�|�8�ȽA�k7�Ӿ[�E!���>�;��38�	8�=�.��.�>���X9-�W�����?���v�t�@��J��4�b�����@5� eU�?�x��Ҋk?�      @/��[W>�                                A�e��@  BL+��  BL��                           ��ׂ��r^�+k�tź��g����@Ai������g�U�yAd��Pe��                                                �_�Q��J��,��/rc��� v��w�#G�ވ�s���
�C?���%޾��HfԪ?���/-�P�ds~*컏>0���g���p�h>�?��$q��=����~��?������,k��7�1?$�����L��'W����ŕ,�                                                                                                                                                �zP�+��r��fc��U��荦˂�@[ZsWAʼ�
7��=Ʉx��%� ��3|>!��L��ƽڑ�d&��<��hh4��� uxy�>5]���ļn���R� ����@>��q[,�轈^��=����~>����o�2                                                                                                                                                ?�w�Z��{f���[�DT>��V&?��U^��ݿ�#5����#+-Z�+�"]�Y�辰��"x�羘��y�¿�+�F���"{+�;C>�� ��ˢ�#Ȼ¡)��"�SӤw>��Zic�u?�U�y����J?��X����I��$����o�&ھ��^�z?��E45�m�I��5�~�a����3@"9)[�  >��x�O  >�RX�����29-2���q���ʾ�^i�[� m���@���ɗ�@-�( �b@�x6� �1���@g�$A��=                                                                                                                                                                                                                                                                                                ?��
`  �"u�Ǻ�>�Ǥe���1`O����U��,�_�H�{�� n1�\8@��N���@-�'��M@�x6SQ(e�1�413�@g��{��@αhI<�?������;M/�l@�ȯ�_j@����aD�?�3�*���A1MTBm�7�[�����j?��������FxAC�r��!	��g$3G�����g۟�'��w'�>�M;K�o�b�(�� [Ӕ��N?*~H�T���ඓr��@2csJ�(@VU�f�X@���hʄ���p}R�@��d����@W" 0U�9?%�2ȷ���%c�@��Y���?�jw�S�)����#l.��8�@����n@��!$�@�P7��A!y��6���WV1��@T]�:(=u�]m�*              @���GMW�>|��U�y@���	| f@��8�%wA��xt   @�8`uR�N@�nr6��@V|�����@�p�T=�h��?xb���?��V�7ϑ�T]     ��ր�`  B��'	¯=@�2�cv�4�G�Z/1��Jp>{���fWأb��E�>�v�?��X�w?        =[�O^HzU?�����?%	W��}佮�Wd������ݥ���ݴ�=�?U�I�?k=��X�t=x��ϬZ4?�����@Y����A�@|����X@�p�z�=�g���?��V�7ϑ?xb���?�      @/��[W>�                                A�e��@  BL+��  BL��                           >Ə���@�r���>�D�њ@����o
<>��=D�o�A*��z<                                                 =�Zq�w @�"d�w#?�߰p9�6���z|Na>Z"���*?E&ƴ���=����촛?����H��&.nFQ�S=�(���=�j�4ھP?%����H��aO?���	�[I�5�1~�>�JXi�>YL��#�ȿ����sJ                                                                                                                                                <�R�"3(>,A����>A8҂bR��3��^<v,\H���=a����<y�1[�>D�����X�<;�����<p��ߎy={x>%i��<��<rھK��s���>�ؤ�@&�����b�.�����ƳR>i �u\��                                                                                                                                                �/8�^aW?>J�1��w���������>��Y��S��t��>xq�ƥR�/8$8�)>J8���>R���L>�:J���.E�I��=���YO�G�-���>&���RE��ʗ���vx�ᡈ�|J��!vM��>r ۊWN�G��,�J>&��~��>>�����@>'�<��|�G�l��>"��@&\�T  >/:<  �}��K�
x���1��o5�T����Ⱦ�x�i@ �﮶  >4��� ?W�ɀBh�?ڸ7��T�5���᷿oU1˅v                                                                                                                                                                                                                                                                                                �H��E~  >?n���� �~(�٪����E�2���� �IYN�����v�J8��� >A��}Q� ?W���?ڸ8��+�5ɢ#���oU�z9@_"�^/阾HG�"��o>~C��y�"@��� #+>�8e�x�>��ZO�@`?�\�ƞ�N��O��/�g��	�W���H��+>AE��??���}%�����d2>0;�.�e)���p���;F�L��C�� �?��<���;��Ҿ��Qd">4	Fq�.�#�Q���?ڸ9�|E��߰M� �o��0�4+�o3�K�5=d��60��=9���G�?�5ң1����;������� �gVK��:�7Bw>!�5~�C�?W��q��g?ڸ3��p�@�Q��׈>@3L��5Bj�gk09<�2�E��              @�GڑPm�sc�7c@���	| f@��8�%wA��xt   @�8`uR�NAa.F�?@V|�����@UTJ!ľ�R,�Aj�?�r�ױV@>���#Zp�j�	���hBi���EO�=d}���и܁����@�Rv��D��shҦ�D��	>��Ô�4�2&?���3��8        =���:�	>F��D�L?L�eڙ_S=��i����:yHg�KOWw�>ݗaU*Ǿc����f>3G#��|N>�oN
^��G5����?��\}��@UTJ!���R,�=�!@>���#Zp?�r�ױV?�      @/��[W>�                                A�e��@  BL+��  BL��                           �)��͡Qe�3
	ud�@����ALr�AnQ'�iN�����E��Ah_�̫��                                                ��|@Xu�C��U�u.пyn��r1���F��������Ѣ?�~ ��=I��	{��{k?�;�H��ӿV���3h`�$��}�E�?25���qn?���Ed,>k5S.&�?�;Q�qB��#��]��?it��~Ͽ�ya��f�?�[                                                                                                                                                �ݫe�iD%���NE�|����ܖ�x˼�f�e7ɹ��I��Y=��W��s�m�WVk�>{XR����זn��l���'����=��X��X�>&�r������b���%Ia��]>�JnBb\����`��>�J�>�C����                                                                                                                                                ?�a?R�g��ܘ߻�l��̟]c�?�J߉E$Ŀ��1�Pω��'�k��
ۀ����Ӧ�kQ>u��<W봿~1s~]��n�����ۍkyb� ���� �p`�����D�|�?�~��c�(�L��m{?�o�)�ԁ�J�P>���q#rc�u��yi�e^�g�5\@��MR�9
?�Ȼ�Lld@d!)�  >��gv   ?a.m]�E���ҕ�鲿{Ն�H���aIϾ���%�@KF,�@kG|R%�@�M�'�@�/�/>h��.Qz�Vz@��W��W                                                                                                                                                                                                                                                                                                ?�����  �pe��f ?aMa�F������om�(�Oʕ/?�Z���0�%̯o�a@kGY�e@�M��@�/�,��.Q�|@�)ᘅ�@ʬ$���_�K���R����`(�P!�@������@��R�I���p0;�OA7�N���������ה�C��%�#cMH�ZAC�G�v����C����b�ө��?��h4	�?����[�?47��	��1��$z1?��Hm�1�������@�.f\�U�@�Tj���vA��S�3��!@��<��@�+�^/1@JɦI�l3?��g�%k��jt֦��@�cmgF�@)��w����N�p�j��1v4a@Y�S9�S��u ����+������,A)"�����G���i@A&�9>8=c�Mxw�              @�Q,6��>4%Z���@���	| f@��8�%wA��xt   @�8`uR�N@�����.@V|�����@[��&=���4���?�?���L?�=� k�@A     ��7��  B���8�@��/O2e@�3�V�
^��?�`Ct���8��֛�Cb�E?��c?��.        =\L��j�?�	�O��Q?%�y�Bܽ���&f���֙.�~D���oF�p�?U�pUx��=���lT6=yI�q5��?�lfo�D@YUےn��@}�F�I@[��3=����"?�=� k�?�?���L?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�+�htsx@�W3���>�C�g�@�(�T%>�l�Ǽd{A�`9*�C                                                =��C�,@Ev�ٯ�?��Y��0W�� %{�>Y���S��?E�����f=�\�
�?�x��6ӿ ��V2�k=�|��&�=�=�e[*?���AC���w��S�?�X�Ά��5�,r>�N2o7x>Y���ou��c�+IR                                                                                                                                                <=p���>+��;�T>`�(�RW�蚪ȑ1�<u�\p�l=b[�_�<y�#�L>DqOH��̽��VrM�;��z�]?j<p>��V�;=|>_���<�ht%���J��s/~�>�ح�^�0���֋t��9Û`>�>i����                                                                                                                                                �-��:��>SOe�+��A�H��\]�ٙƾ�W.`���>w�Q^���-�dZO�>R�NN�>Q�����>�]�ܯ���,�L�eG=�a虤�FGF�.�>'.�m@j���:�T�D'����V%#��~#��T�>q\š]e�FA��a>'.��ძ>
q���>%�*��8J�Fv{Q� >"v��!�@&\v�  >/g�m  �~����������v`�U�~�b2��ђP��@ �;   >4F��  ?W��A]�P?�p�����4+�TEAJ�n#�T�o                                                                                                                                                                                                                                                                                                �Glx0�  >?���@ �~����zT��+3j�)��r��նA����2(��H��_  >Bzpߠ ?W�ҬnA�?�p�߹C�4+��X���n#�օ�@]��X�H�Hf�� 6
>4o����@����y*>Л V���>�A�Φ`@_*(/J�z�N��s���g��'�˿�p�	��AD+�2�h�?��uRF̢���Y�v�>0KƴH����`/�2o��<I�tܾ�r���?�<���^T���\D��q�>4)�M���#ܣ�:-6?�p��]&���̓}5׀�n��.�]^�m��j�$�=_)G�T��=2�сP�?�*G�C��t9�Qy�����~����g�>"M�>S��?W�����?�p�u�B@9�e�>@u�FE�@_� ��� =�[���+�              @���M�:>��L0��/@���	| f@��8�%wA��xt   @�8`uR�N@��L#A
�@V|�����@�r��=a=��ap[C?X�5&?�њc@��@_�     ��p��   B�A�po��@ե��=��2��'����
܊:	��_�ZV��Ab���	�?��m!�;?        =\��s8�?�<�T��?&�s�`�x��̹��@���.��<��`�Ub�?U����=��`��3�=yԷ�hR�?�͓f��&@X���P@#��4@�r��r*=�k�׍\?�њc@��?X�5&?�      @/��[W>�                                A�e��@  BL+��  BL��                           >��6�T{@�	C��`>�HϏ�G)@���*)��>��l�(�A�ŤN��                                                =�W_@��J�?���8����8�>Y@�.]�?F���U�=���nM�?�Ћ�$dd���^ xH=�"@w��=���ZM[?8.�g���'�aXp?�� �:fF�5�V[�%>���H(L>Z���t���0)Q�                                                                                                                                                <�qz�:�>*��>>���o�c�螸T�><ul�.�=bÞ�b	�<�yX>,�>D9�tx���Ѵ�;|^M���c<o�����=|�Z�%��<���QO��Jb%���>�ضU�,���_����Ѱ6��K%>jF�I{C                                                                                                                                                �,�A[	�>^�������X�#фN��R8�6
��o��[>v��1���,�����>^>>P���}<�>���_�X��+�Ə`��=�Y����E$Q߷q>'`3[0)����ˬ�i8��u�U$���>f�Q>p��ǻ���E$
=��>'`'���,>��Xp�>$��>���E#N�]�I>"�n�#h&@&\�  >/�][� ��D����h:ŷ�WW���ѫ��ْ3@ ���  >4z��  ?W=��7]�?�/��ؑ��3V@6X���mC��                                                                                                                                                                                                                                                                                                �F1���  >?�o?@ ���� sr��nI�NM����	����r�d�G���0� >BAH}H@ ?W=�9��?�/�ވ��3VwJ���m�
�@\�9)�_X�H�yx��l>�!$|��@�z��>�
���k�>Ϛ77�:@]�zY倧�O/����g=��3���/�u���ACVx�Q��?���~�}��7ف�T�>0]]�ʽ�!��^=J�<ǅ'(�����	���<l��s�Q�����ƪLl>4L/��vY�#��S�?�/�؝����!����m�ˏYNm�l�D�+=a�z4oR=K!`Rh�?���Eצ�����u#��kW��I��c��>"��_U��?W=��FR?�/�6?��@FH���G>@�&�?@h����=�,#��]              @��Խ��>�1���@���	| f@��8�%wA��xt   @�8`uR�N@���9��@V|�����@D%,?��=�^���a�?�4}��?�f�q��@h�    ��^�v  B��V6�)�@�Ÿ*��1��.�|������ޮ��1����:�?Fe�d��?��vLU[�        =] +eX�?�wFWm�??'���`���ѨҹE�ב����"��ح��?Ue��Ś�=��9�%�=z`&����?�5�ѣ��@X}Z��)7@��k�n�@D%,@8�=�^c�W^?�f�q��?�4}��?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�s��5ư@��Lb��>�TL��@�[WZUY>���s(�AJ�xջj                                                =�`"z�9�@"Jځv�?����Eʽ��}��>X�[�(��?F�f��"f=��gZ?�0zJc�-�~�%/"= D�L;b=�C��eEf?��ߗk}��=�v�?�z�hO�\�5�-���>�lQ�/>[d�N�i���@^�7�                                                                                                                                                <��k5?x>*j����>��ǻ�g���<u�{=c+�ӦW<d��+�>C�$�7���Q���B;t���|	�<o��M=}X�)�O<z���Q�I���0w>�ؾ��^���G���(E�:,>j�(�)j�                                                                                                                                                �+b�.�>k���Ľ� ���4��+S�:���YNM�>u�����+b0��s>kVu�.>OY��2CI>�L�A�#�*�]BY=�^	ȯ�`�DJ�f�޿>'�b��P��ɑ��>  ��)�\�5Z��[R��>p)�5��	�DJ�D�%>'�V���=>:���{X>#�C~�<�DI޳�.>#3�㗩�@&\h�  >/��͌  ��h՜��(���Hhn�$�XEwV� ���{=�C@ �.�*  >4����� ?V��Nm#?��8��V�2�V��9�l ���                                                                                                                                                                                                                                                                                                �E.o  >@O�  ��s�����@��}���Y�_1��.�={�|�Ft�hx  >Bj{�O` ?V�0C�?��9����2��s����l ,�@[^��b�H�~R��>���:���@�����7�>�����>�񰉃�2@\�ӏK̾Ox�����f�4�U���J���fAB���aQ!?�*X㙁�TQ�o�>0oe�u! ��[��x�T�=���=���Y�l/��fE�侢.�=��>4pdU���#�==��~?��:��u���j���d@�l�DBtΊ�k�ʎ/�=Y1��r�T=5J\�J��?�{m�脾��R���,��.�D�\s��I�/�>#:(�
r?V�+0��?��3��u�@��Ex�>A��.�BT�@[R`=�O?�3&              @�"F����2����@���	| f@��8�%wA��xt   @�8`uR�N@�1��ф�@V|�����@�����%�!Aqw�?�f2_�@#x���A��E���.�@BQ|��y�E�a��7?Dݨ���wD�����6D��Eb1�YDu�~L��C�Gӵ�N?���3�ӗ        =��$x��>�6q� �?L���%�f�ӑ���D&<��ol� �uv/\5�>��5J2�{>`�/���Z��
:@ ?��?�p��`��yM��^�i� F@�������!Aq=9�@#x���A�?�f2_�?�      @/��[W>�                                A�e��@  BL+��  BL��                           ��{��B��R/�+�?�@��'�O�0Ae\,u��@7/�]*�AVFc\�$                                                �Q�ͦ����-��E��3��q�����ʷı�>�۰L��?�Ͳ��Z>�rl�4�?��/���9�����R�����i�E��zx��'�?���籀p>��h�r?��_~�3_PV����X�Ӆ?!/����^����                                                                                                                                                �nM�j�/��Aɂ;���#��u���G�U=T��JH�=�I ,�=t'����>2��Μ����wJmgE�7ZVպۣ��1��M��>E��K̀�/��t�%%�Ix�>��E���=="��� ���E�4�T>�R�I6                                                                                                                                                @ Jx^�m2J��~��
$g
?�]�]��ſɅ�!��l?��EMF���COBC@�uq�z�8���v����t��5���y��f��u��͚�e�2�ɳ��y?v��e?�	�= �S�?��l�B��uV�����p�s��DJ#��E�X�u�/�߿�X���?�?��Zq��C�G�V)?��,�;��@%m��   >��|   ?�l���T����	FIv{�Qb��`T�M �������"��0���v���z��D)@�&�/�5�1�iCS��I@C�:�_                                                                                                                                                                                                                                                                                                ?��R   ?_�y� ?�I� �����Yڅi��B��	�\��s��u����$��m0��ou�Ƹ��`33��@�&�<��1�]���H���GV�@�#�/�@ʜ�;�#��(>��~�@�%�7��Ӏ$&�4���e��P�A0�K\��@�)������
3��^���ӢcZ0AAb���<@�hB(@1q�+ƫ@(�nyԠֿ�QdW�?�VQ5�:�"����e��$r�ic�����C{���?�˓pD��@���c�@Ѣ�������X}�9y�0���@pv���ke?��}÷�P��R0����@���P��K^+&E��#e����.���ց�S�$��R�[��M�D�@�u����@�m��y.@0�C���&@Q@��=w[]9�;�              @���|?>�J
��{@���	| f@��8�%wA��xt   @�8`uR�N@���y��@V|�����@��h�j=�-��(O?�D��ݎ?��lΛ���Q@    ?�{�mh  B�r�]�`5@���%�t�1&�.	���Cq��_ͬ��<5�L�]?��~ϼʭ        =]|_E��?���Wr�R?(�#ix�����>�Eŭ��qE�j��V��v�J?UI����=���9Y/=z��Q��?���f{G@X�q3X�@��u�M+5@��h�H�=�.#���?��lΛ��?�D��ݎ?�      @/��[W>�                                A�e��@  BL+��  BL��                           >��S��8@�{�jr�>�2�n+nA@�����;T>�|Ɍ��EA�q���                                                =��ڲx k@{����?�)�џ�����bF>Xz��[�?G��2=��<����?͗�g���K�*9�<�~đ�c	=��=j�
�?yP����̤�s6�?�4�__�5�����>-��� �>\p���4���*�}�?                                                                                                                                                <^����>)ܮ'/�j>��~kN�谛����<tĢ/To=c��uK_�<�똲>C9�U�̽l�I_r�;m9a��w&<oy�v�.=}���^J<9Ls��վIJ��p>���?4����Y��2��ҡ�e�'>kh��n�!                                                                                                                                                �*G�)Z��>{�2����ec���w��Q羨�i��>u���P��*GNw#6>z}=+��>M�T��k�>����A�N�)v��u>�=�Mn�]��Cxgk>'�."�G[��DՕ��*��x6�
�����Ca�T>o?T�-���Csh�W�>'�!�v�r>�� xR>"ܔ���C~����[>#�ú~��@&\��  >/���  ���u�[��=��3�Y�rբA���̅�u@ ���  >4��@ ?V��/E"?��y{n�1՘sF�t�k
%c                                                                                                                                                                                                                                                                                                �C�`�f  >@��  ���k(�]l��C,�[����f����O�E���EgSJi� >B�!�� ?V��B��?��zM��1��,9+�k
��,@ZH;D�H��:�4>�!f�@�NO�n�>�S��>�$�4�!@[��]���O�<E���f��^�����/�4AA�̃�0,?�r;��+��
㍗�&�>0��[�!��n�iH�>eّ���f�9�<���������g�o��>4�^�;H�#�r�'�?��{H�8p��̕���k��g��[�j��*\k=Wwz]��=�̖�� ?��`�#���K�]�(��O���:�ҁhJ4�>#�
5�(�?V���c6V?��t�!2@��n>AK�+:�HA��E%<�ŧ:V��              @�w!�\���6^MG@���	| f@��8�%wA��xt   @�8`uR�NA��8Oj@V|�����@3=p�!�`,��>�?�+^��@)�[SF�
��%?/� ��c� |�E|��DQ&NX�D�� ��4D�ba�"�D|��F7(C/���i�?���3�b�        ��FH�>��>���?L�$���T�e��<3<ߙ���Z]�m���a)>��Q�+�?=���PAM���R�2�?� �j(*�f�:Ƹ�����ћ�@3=p�!�`,�΍�d@)�[SF�
?�+^��?�      @/��[W>�                                A�e��@  BL+��  BL��                           ��W�#���VԑO�@&Yc� Ak;8Xn��@%W��Q��A\�XjN��                                                ����읋�&��^�H����ٸ�7�CD�R�FG����u�?�qw����>wՈ��?�EpJ���s���}�'Z����`���c����?�N
�*�=�����[?���!����2<�6�E��T՘�?Kʏ���lQ~c�                                                                                                                                                ����K�5���{�����@9yw�y�`X��	����V���n�=�H{J~;<����Б�>2].��;��HT�g��W+����6�}�"�>�K׼/�m �嚣�$����>�-@H�"�=�X�������pR):>�� <<��                                                                                                                                                @���F款��Q�[��`\k�gV�?�K�ҥ��}r�b\��):Q>��@Pl��T�����
��m�������r�?�@�t!{a`>�V\{�n�2:�L�Lx>�(8$�������?�)�@��~M�r�%�5���׏�D��gby>�< aҾվ���Ӎ�?���3���C�>R?L��	�2@$ăD  >�F:�� >�[i�u8��ы�߭��]9'��K�R6*k�\����%kX����z?�����§ׄ�@ڼ�BW��/� �:o?�0�U��?=                                                                                                                                                                                                                                                                                                ?��@  >���\� >�'5�������1)}�q�W�O�W�m�8��迸��ŤV�����sV��@ڼ�����/�a�W��0� ��@��P��?�0��ʿ�oU�fp�@���D�y��EfCK6����Mk,AIK�ϼ?֨�p�@ TiD�)f��W����A@Ly
jm�@e�z�qe@��,�z�?Z��/2
$�	V^��-M?�[YW���׫�g+�n���s����G$;E��Qkd������H@�	=r�o��Rք��a
�-�wV@dP�5�?����	��f{D��@�GLq�W�.ͲYxg�d�e��l%�KU �����4ln�H���j�kx@�Ԝ�ϟ�A2�{��@	a�-!:�@bv=�~=����ZВ              @�o�ɂZ>��_���@���	| f@��8�%wA��xt   @�8`uR�N@��p[�r@V|�����@(Ɏ�Z'=�{�]�?n�D�?��r2���bv    �� wĀ  B��Uq��0@Х��ٍ��0z���'����������~�Y�9��>?��?�����+        =]᫷@�y?�Tt�r9?)�pED9��b �C���؟V�'Y����_�,o?U-��9Zk=��L#�={����?�`ޑb_@W���:5�@�A��0n�@(Ɏ��=��I��?��r2��?n�D�?�      @/��[W>�                                A�e��@  BL+��  BL��                           >��T�W�A@�<H�f>྾�;��@��(��Wr>�7��ܫA ʎ��ݬ                                                =�J�Ӂ@�@J�*?�bѝ����)rՙ$+>X �\�'v?G����=� ��n�?��K�{>�!'�)�;<�MM�=���D4�?�ev�ὧj�dZ�?ұ��K�q�5���.>g\z�>\�r��>����x_f                                                                                                                                                <�Q�P3j>)VO���> r��\����	��<tx���y�=c�e��z<��(��l>Bژ©��=Z&��i|6;^ ׆�҂<n�� sug=~�����<$ ';H�}FcN2>�����p���)�s�ϼ�=���>k��&ݏ                                                                                                                                                �)?��{ �>�mp�x��bq@����r7�d>о���n�>t[<`{_�)?� O��>��w�6>L!O����>��Ee��(~��TS�=�!�^�NR�B��+>'��o������!�ܿ��ͩ<Ɏ��b'�k�>n>6*Z���B��O�>'���W�:>��5rt>"��D`��B���ķ>#�Rl���@&\_�  >0��� ��a�%�\����jgG�Z摡p�׾���}f0@ ����  >5"Ȭ� ?VI�nm��?ّi����1'����j$z�w�                                                                                                                                                                                                                                                                                                �B����  >@9�K�� ��l�(ߞ<���N�)=��N��7ON��o�����Dk��� >B��~<� ?VI�&>`l?ّj_�kn�1( _4rѿj$yA �@YD  zݾH���w�>���f�
@�A�Wk>�6/	��>�O *7@Z�b"m��P
xׅ���fI��,s���|Z��AA(!�>��?��o$8�^�	�;=\;�>0�?�'1�q��a�p�??���\ʾ�N��«<�n���~���6mY�>4��ax�#��L�j?ّk\�����:ZJA��j��_q��j!��L��=RY�-�9=h{!�� ?��ݧ䳾�Qa�X���o�' �N[�>$;Q�Lc}?VI��L}S?ّc���i@���>>A�L��BGx�fPG=kR��K              @����fQp>�w�?@���	| f@��8�%wA��xt   @�8`uR�NA����|@V|�����@��h>W3@]��?�H�s_�u@/��q��Gv���`A��d���@E&�4�c�ȕ�UɦĔI�����=^��D�NL��nCFk��=�?���3��x        �"h��>t..m���?L�@�ZO�sm�YS/E=�XM>���f�\|�C>�w�\d>q5�8^����{�?	c��`��a����n�?u��fq@��h�>W3@6E��@/��q�?�H�s_�u?�      @/��[W>�                                A�e��@  BL+��  BL��                           �	*��ș �a�NӋ6�@B������Ar;�89@Ac�7Q�Aa��s�                                                ���@v����:l���?����X�o�f�<6>�])��?�np�<�>�A:4�b�?�j=Z��h~�Q���2�5FQna>�4ٿ��w?�����ԩ�|gG�?��A΃��0�9��ݾ�޼����?0o+i��\�B�                                                                                                                                                ��xF?J�t�#����=�#v2~;㼋#��E�=��2Ԧ=�ᒭ��H=�l��9>4g��|����R"ʗ���Z]?�=$EE���'>u?�F(�<d=��S��$�?S�q>����m�=T_�@������1�>��m��                                                                                                                                                @#/C43c\�̙��6y��1�8�N6�ӛo��,ƿ�v�As3�?P�Gh@6��B�0����n"�����yq&�@忺���~@7X�>�.�ZX8f����3��t/g�?��EKپ���c� 
?���X?TP�d{SF�?#˺��D,H;}�x>�#(�C�b>���i�[?���gԌ�DY�Tz��BSK��@$���  >���"� ��7��#o ���'޶���e�sKOϿU'Χ?�t�cNꋠ���#'�=���0s�@����,k�-g.�mԻ�F�,�9�]                                                                                                                                                                                                                                                                                                ?��D��  ?S�Jj� �� �gC�Z�����8�)��.�ٝ�QYNE+]��v\p���P�����0��>�N@�������-gN!�q�F�s޷�@�L��A��w1���?*5��kG@���L'&O���N��?����"A y���0D?�ITN��@3��?�U|��1���A>�y�pf@p��VJ?�����K�;��Ĥ>��
��6?y�~��+���j�*?<v>�
����L(ì���@����� �Y)扺@�&q�����Qh3�e��;�Z@Z��;7?e�4qp>׾��0�8@�5���^�9~����LD(H�>/���'���N�8�a���4E(@������Az���|@)�]6&}�BƘ���=:�~y&*�              @�����|���.��^�@���	| f@��8�%wA��xt   @�8`uR�N@�P�[��T@V|�����@���چ��#����^?~_�(���@ ��*@a����� Bz47xD��D����<�%{ ,Gđ���K�Cwo�m;v�P���LtB��E-���?���3�G�        =R��2�>�Y|q���?L���?��=B%��q=B�� �*v$�x�n{�->�����R�ȃ.�4=�Vj0�i|?~<��R2?��ey�?�\�A��@���چh�# R��8�@ ��*@a�?~_�(���?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?�2V�
j�q��hJ�Z��� ���Aw	4��@��oA�O�CAS��v3A                                                >��u�� )�%�#yz8��ѨU������˘}m����On萀d?��^�?��R��K"?�{�!�c�?p0ǒeY����G�>u �g��?;i��X�=�����:?������3�5�}�>��ik���i��|v� ���6                                                                                                                                                <�6s���ԾBX�/����3N�׼2E���+�*��_>ɼ�)���}��3`�>HV��=��D�I��K�>P'<�I,.&�=��s=�F�1��a�A�&=���q>�+�!�1�-Ӭuϱ=W��msq�>�*��B�                                                                                                                                                @A۞(f�J>�P2=�宾!��ak�?�)@�n
�}^#���ʒE@8��\x�>����5���3���]?X��b �@9`��ϣ?��m���G_��־�QE�s>�I��[�+8��x��3 ���EJ��|)>ꎄ��M�Cw�2�MӾ�H9y�u$>�5X��O�?a��ǂv��Cvp�8������W��>@%����  >����( >�skw����c�=V:�J�l���f�H��_�,������{�?xV����?�>��f-W@ǉ%�g���/�Kᭈ�@�Mr�8�                                                                                                                                                                                                                                                                                                ?�u��@  ����E� >�7��	��cH�P���� �Լ��I�X|������S��X?xU���?�>�[�@ǉ&h�	�/�d�	G@�r��-@��X�F��:��~J�}�R��Y�c@����=
�sĢ��U�V�2�tkA����x��zh�:��㲫������+&�4A@�p�����D_4ܤ?�
?:�K�>�c��D/�=ʏ�-��?E%B9m�1N�(��>�}G�Y���ݛ��X?}�,	xV�?�� �ƛ{@�����Se����B�rN@m�)(���V?*��<.>�a}��tO����`�@y�4���?��E�Ze�EV���.�.�*��?�V�"N?�CD��F�@�x��ͅ"@���`�.��(�JƠA�|RotA2=6/�?�
              @��.��m1���1D6L@@���	| f@��8�%wA��xt   @�8`uR�N@��ud]T@V|�����@���ľ���68�?h�G/�@���e=+A�|?^�@ AM�$q#�DV�G� �B�Zl��V�fyĲ�C���DVb���rBoh6\[?���3�u�        =*�ӏ��>�\��C?L��,��Pl�����0��|����0⠔?N���]=�D���=�O
2SI?1��)O��NT'�֊?�U�%Q�@���Ѿ��%#�&@���e=+?h�G/�?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?���Y� �T���%<�_B�,9A]��E�;�?�Y�G��A@����4�                                                >~"9`�)-�G�̲'p�Pf�����fLo�*����p����?��ZC�)������?�_��+Nj?d�#M��Y=f�Z�m�I>[@}�y��?*:��m�=�E�S�<?�?(5�΅�4�F�7��>�$����i>��t�z�����̠7                                                                                                                                                <���_��v�:��|dM�-`�~<�����?�?_��^���	=�a!A�Ϟ�*z�nz�>C�B�=ڱ�Œ\�;�ϊʠG~<ѳ�N�܏=�	�p�e��)���ٿ	�&��j�G>��ndxr��9^I7H�;�4В��>���`�                                                                                                                                                @9�J��>��������k�?�@,��=�D��)
�듾��Q�9e�	�l���>z$ED����q��?Œ_+o�u�!�Ǵ�����to�LY�B�ؙ𼥾Qi���%=�q�,������~�U�G�y�@�>�:~@#���B(F<dS��P�[�~��>h~�B��>�y�A���B'�E�\۾k�D6�@&= :�  >�f̫<` >�0g3:����&?�ÿ"zG����4���yXF��@6�]  ?8w��?�ĺ��J@�i�U�9�0UM��O���cy��                                                                                                                                                                                                                                                                                                ?��`  >��(�l >�>�������R"��N��7%m�v��5u3
���SzAZ��?8x�,y|F?��Q����@�iᠥ$��0Ux��$��c���@�] ��l?ߺ��p���ڋ7LNl@�������O\�n�6*�Q� wI�@� �| >i�RG��2��� _F"
���X��.�A@]7��ڀ��3�Q�*?��V<oX>��v���m���s���?�c��2�d��TB_������"M�0������?9so�'�?:�W�0�@�wav�����ݒ���f?Ԃ�� �@\�]}*2+>��$�#/0��+�~��@W�`�-R��
�1�<�89g�q	����ͅX�?H0@���?�9�̿U�@��$'@�\*0��?ZK(
T;@P���y�=y��rZ              @��c�6>�V�r�'@@���	| f@��8�%wA��xt   @�8`uR�N@��b�@V|�����@�ԋ�
=�y��9�?������?�O�6��P��    �̴��h  B��|��@�,����/}��+L���gc/�D��;N�6�.UGb:?����d        =^C��,�?�3�iS��?+.��#���5U;�=���3"c�:��I�,�h?U
dϿ�=�#g���=|3[�w�?�w3��Z�@W���lj@��u�W��@�ԋ��=�x�ޏ�(?�O�6�?������?�      @/��[W>�                                A�e��@  BL+��  BL��                           >ʭ�Vd@��1%O�>�lY*G��@�C_���>�ǧ��A ��/��                                                =��eϗe�@(&�T�?ℝ������B��@�>W�.5K�?H�P2k>=����
�?�_��S_�?*?��^ܼ�N���>�=�@D�=I%?_�7\,��9@��B?�Aq��G��5�+��>��	&>]��?I̿���N��                                                                                                                                                <>m��>(��'�+K=�k�d����*g��$<t#k�-�=dtbz���<�z�Ϫ0>Bn0q��=~(/n��@p]��Z�<n4����=PX�P< Q�o�H3P@��>���G���,3�L�
�Ӵe���>l����                                                                                                                                                �(]IK>��g?ɽ���R � F:������VcT.�>s���=���(��|L>��̬��>Jp���э>�k-�����'h��=�=����A�>@"�>(7��j�ȫ�C����5��k���)TM;�>mS2�6�A�9�z0>(7���	>�vB>'�>!e�l���A�ey>$F�8!��@&\��  >030�w@ ���i.2&�����ى1�\��K�u�� �Ay<d@ VU�  >5k�"�� ?U��ϓ��?�_�<-s�0d���>ƿi#R�둻                                                                                                                                                                                                                                                                                                �A�OT�  >@[�,�� �����-��b&,��q���Su�јH���CRa�  >B���̀ ?U�Υ0��?�_������0d�Xiſi#Q��@X SQJᑾI"Yn���>��w]h,@�"!]��>�=��yH>Ђ�6͵8@Y�F#��P=��w�e�ʴ�[Z��_ߎ
DA@d����5?�
mDk:���E�� >0�J�2&i=uU��*��@(j7(��q��۴<���m8�����[�o�>4����X��#����?�_���<�����8�'�iѓ�X���i5.�bi=d��-��=^4�Dgd?�6�v�\���t�8ٍ%�јA	��+�tL�!>$�y���?U���h�?�_�+�֜@q#��T�>A�{�}(B?� �D�<�aA`c�              @� �)�Y���ݫ�ɓu@���	| f@��8�%wA��xt   @�8`uR�NA��w�@V|�����@"F���(�=f��[q?��syp�@7o�3�6v���M� �>�E~qoE+��$_�_���ޔ;��E�y�D�c��=\D����<���>��'�Y?���3�@�        =p��
{)>]Vt�$�?L�\��!�=���qw��=p4G�]�W�0v5?�>�`�T��xN	������}|>��'�33�XS�K6b?�cG't�@"F���'�=f��]P@7o�3�6v?��syp�?�      @/��[W>�                                A�e��@  BL+��  BL��                           A7�W��Aa��ՙ!�7��W��AMk;G�~�@Pp��<FAfSf}v#�                                                ?�_e��3x@ Ý���g
��?����hD�@�4�@���'��|^,�[?�k�
�\��bƥ���?�:��4�?(�v<-?��?{��M>�7ƙB?���;j�F�*��]�5M��9�җ���м�d#����hl                                                                                                                                                =�!�ϵ�>:��f����H�=�q�&u>���^jj>'UT�n�ڽ�;[� ��>���-��dtOp�]={�~��(=�OtcGN�>Yx{PĽF�of�{e�"�]�&z>���ȩ�C=mv\�O =F0뎁�>��m��                                                                                                                                                ��/o�?�1�Um�<?��Y�5�+?����h���&%�̗T�@'�ޞ�}�N3�4��@ gY�Bf��zB��W��'4s���Q�,��_@H�Ӽ����]nͥȿ�g�6u5?y���l?�H���#��7�9�W?��&���A���N������R�?(-��
ˣ?����ahv�A��K۾����zJ�@!�x�  >�n�   ?���B����a��J�,�s��)GN�["�
<]��������PW�~W� �k��/�@�1m�`�)*SL�N��MJ�l�.�                                                                                                                                                                                                                                                                                                ?����  ���P)� ?ι�����_���Y��1�g'i_@DWԦ��c����L�rd)���" ��+?@���"�)+'���$dLh�@��H��9����+�� �T����?�@�O��@��#p������7�� �A+���J����� (�O@�+�{_
�'�WR1A;d P�n���߭ێ���!BQ�@"Լ�?��$/�ʈ?����E��]���Q�@:��}���A����@G��i`�
@J-=\��H@�f<���2�55Es�5@���)1Ǩ@V���\�0���f��t�Uv�@���P�On@3�K�q*[�,,Kŉ2��4?�yΕ�SIw!�<$?�̳9�@�ǿ'x�cA����(n�%�� �6�@X݀3mL=���}�              @��/ї>��%�*�@���	| f@��8�%wA��xt   @�8`uR�N@�3�!�ש@V|�����@!d���=�ǎ�w�?D���?���OZ�X݀    ��I  B�?��+@���Qm��.czS���N�^C����嚓N\�4�����?���Xb9�        =^��zC?��~|��?,8(��0���2ђ�ٰ���;���v���?T�����=�,�!KW=|��$?��A�|�@V��ɿ��@������@!d�n=��oF���?���OZ?D���?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�kT(���@��&?g=>� �}q1�@���n�r>��Bs�v�A N<8A�                                                =�X�]��x@��5�L?��Qy@ƽ�\��<�_>Wn�$+'�?H�U�!�=�*��˅�?���
<��?�Tcp���ڞm{��=��l:�[�?��\_M���D��{�?�賅HU�5�mˮ�>9-H�^�>^z�|��׿����G�                                                                                                                                                <��mŝ�>(C���v=�IP�ֻ�����<s�1B��=d٢�`��<2�<Rr�>B�H��2=� |��-�cd_�Y��<mع����=�*Q�(4< |[�?ٞ�G����UP>����d����\��_���3��K�>m2����                                                                                                                                                �'4��HD>��5n�"���z��d����/ཋ޾��z�s:�>r��q =�'4��T>�����4>I)�$F�>�j.���8�&��T��=������AGb���w>(m��8�t��m�L����8���w�OQ>l@��"�+�AG^^?W>(m���v>�Ac~'> aE�dXq�AF�Q�;^>$�\A�F�@&\t�  >0M�@ ��{���t����IG�;�^$�� ���>��R}�@ k�7  >5���� ?U�c�Ì\?�<d��g�/�`�{�h]K����                                                                                                                                                                                                                                                                                                �@�|9�� >@y1��  ��� {��Z���x�܀澫ˤ�b�ѺIjtk�Byg��� >C'o�� ?U�qm%
?�<e`Q?��/�k�r�h]J8�@W?-pMU�IKy��܀>��#��9�@�����`>ˀӑP�p>Э��~�@X���6��Ph���U��e�k�=H��<xx݌\A?�m�7�G?�q��g4��+��Un>0�;�-=���2wо@���Ojؾ�ˤ��Q�<��P.؞���+�Za�?>5cl�P��#��eA�?�<fa3+ƿ�7㹰ؿi�&��h������=ec���=_��n)�?�7ͩ�kѾ��W�[@��ѺB�������Z��>%s=9���?U�k�=N?�<^D'�@��r��>BN�oz�ABb�Fi�*<����] R              @�um�A�Y�I{��@���	| f@��8�%wA��xt   @�8`uR�NA�D�]�@V|�����@����Z���/fh��?��2����@<�bm��kBb�Ǉ��R�0��QFQ�E7l]��7�9w&,�#��uA.�DH���Z<D�����nux2�T!?���3�ʞ        =B���+>O:,�`�G?L�d�5H=v�n���A�I>��6�Nᑫ��)>�@�VRl�^W'��=����²>�GeΫ��O"²�?�PkK~�@����Z���/fnl�@<�bm��k?��2����?�      @/��[W>�                                A�e��@  BL+��  BL��                           �5U{��rJe���k6.�&OAl�y(F.p�k�ck>Ah��]yt                                                ��5��̿��sMɖ���)���;�a�9�Rd��ڊ��p�s?��r\�����ϙ�!��?�՟��W���MTR> �P>>��xՏH?� �[3L>�l�)M?�w����%!D��?co��30�M�shp�}����9�                                                                                                                                                ��}MQ:�V��oK9o"���h�3�
�~l��¼����Z�=�ǁOT^Ƚ!jY�T,�>"<O�T�t�ν�D<70<�Ӏ�0^q=R�{��>�> ������V��پ �p�4�>�m����*G�(��=Ú��u�>��XB&�                                                                                                                                                ?�pi⍦ ���uv�p�|��١��?�Σ��oA����t�ތ���
���!�!;G���ʁ�t�>�Xb�u��Lh�^���"sɗ��A�����!ߗ�ښ� uwE^�R>�=��ULm?�ɥ�B3,�}�1��?Q�Ƈ�s��C��&�C���(1��>�/��«?�1ZW���D2��?mHu��~�@�%t8  >�B���  ?������?�Z2��zY��2��]b�.+�� �j:��@����^<@0�޴�@񈖅.���& ���n�@d���hV                                                                                                                                                                                                                                                                                                ?�L�   � o�I6� ?�A������>��u��� hc&r��HZ��v��n0�@��h`��@0�l�N@�h�W�&����@d�)o��@Ɇ<�u9�ˢ��Cx?=��:�X@����ڢ�@�1���s������A0N�Zki~�C��z(R�l]��J���E6A9Wa�T�����jk�J����7�j?L�6�����=1ݪ�i[*;�d"�#Y?`ITM?lZ`�N�J��0"� y�@=��;�i�@X!Ȱ|@������	W��U�s@������@LbKl�p�?)��d����*}C=�@�^k/�U�@<-[�T�8��L�W{=�A@2����z���-��_��t�pA �i��E�_��Wx@_�`o��=��X��9�              @�n��~�>�[Ks��@���	| f@��8�%wA��xt   @�8`uR�N@�RK�ļ�@V|�����@����i=��=Ŕ�?Ѐ(8C�?�����vy@_�`    ?�0�  B��vt�@��V3݁�-a+K��G�����������U��2à�߮o?����2��        =^ѳ�-ʏ?��r�w�K?-DG6�H4���i0Z��!(��K��i���X?T�7�Q@)=�5�И�=}=�<ϔ�?�|M��J�@V;���c�@�D��y�@����"=��t��ݝ?�����vy?Ѐ(8C�?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�/nm�[�@�����>��8�0@�����t>��`/�A FE��                                                =�ظ11��@%���V?�8��7y��y�j�w�>W%��7k?I	�c%?=��Z�b�2?�^;���)?{r'����O��=���2,�?	�,6Ƚ��&��P?ѓ�sa��5�a��>��O�>_=�N���p�,�^x                                                                                                                                                <�|��>'���2,�=�9-�;��������<s����N�=e>^<�>�� �>A����=�P\�]f��r�f�F�<m���jJ�=�B|�!)�< �:]���GMN�&�o>���)�����髪n{i�Դ�"im>m�h�0�i                                                                                                                                                �&_)��fb>�$]q���A���&E�"���0��G>rh�*��&^�,F$:>̈2��w>G��|��>�~x�|,��%��e�T=���(���@���B�>(�_��ܽ�4.�l6�չ��!k���V �>kq�w���@��c��>(�Q�oe�>�Ų��B>wC���z�@�@"H�>$뀇�1@&\�2  >0iIy�@ ������m���ːZ�_����6��]T���#@ W��  >5���� ?UsA�[�?��j��.�*30�g�gg9h                                                                                                                                                                                                                                                                                                �@-}��  >@�ad  ��Ѭ�U#��"4a(+���3g�r�~���͑�@~�A�k?#� >CX}�*` ?UsNhl��?��أ��.����
�g�ߝ�@Vl/�[L��Iv'ٯg>�s��e@�*斋gw>����|&l>�י�iW�@W���VF��P����3Y�esFHeKw��b��2A>��H`2�?��a�N���dCSA�>0ߵ�{��=�B���i��A���i ��3g��e�<�ĉ��ж���R.ȷ#>5J*�X�#��
C�U?�	�����㩨�Z`V�hU���@G�g�IH���=`[�y�J=Y�]?/x?�<CR~+���6�q�����ƃ3v���I�U>&	녝�%?UsH�v?�S���@І���>B�Q�ӗ�B���4W�=(��f]�              @��j��� ��y�VFG@���	| f@��8�%wA��xt   @�8`uR�NA����@V|�����@��7�9�Jv	B��?�o� ^2@E�UC��B��`����R���T$=EZ��?d��8Ԯ�[.�,l�}��%E+J﹯[%D���IjF����]�-�#?���3�a        =�8�@kL�>*��ռ�#?L�lK�v�=�F������8E��w�3�F�7\_>�?^��(9��!گsg�>]��!>��h�UC:�5��'��	?��K����@��7�ٿJv	>]�@E�UC��?�o� ^2?�      @/��[W>�                                A�e��@  BL+��  BL��                           ���r ���)�$0�'���Z�+%('Ap7?s�^����#Ai��Ws�                                                �%�ɍ*�׿�!��P�v�k��*����f������a?�&�V ��&h}E��?�~�TB�I���쾃Q�G��?�Y7�s�?�Q�j��>��d�0ң?�<��&��6�YS8?��#r5ޑ�ƞ�G��U�
 &#�V�                                                                                                                                                �B��O���+��W�b�����G����܀.ν:�eQ��=��_�|��p�>��ea���H���Z��5J:t>ts�>2e5(?qu�I��sK�,ǀ8�>��!~������'�>=�gf^�e>�;Ռ�&                                                                                                                                                ?�_��w{`�?�������Ը3
?�Z����r��@�8�<W�g��P�Q�pF��;s�
�>��lI�d�y���LE���mJ����0q������f�d���k�tq�Ty��Y^?���q���0�5���#@Tkˉ���D�!ɮ�����=mȴ�{-�ϰ���,���S.�K�;�Ͽ�@,�3U�@5ď�  >���0   ?�")G�"���G�u���X6�;��^qpf-3� �^��@�9)G�[�@� �y��@����½��!�ǽ�D@��N��9                                                                                                                                                                                                                                                                                                ?�1P�  �����	  ?���9����F�4@��0��uNQ�@O�K�1��  J��@�9u]�@� ���@���)Ri~�!�:'��@����P�h@�Jr���@ �ݽ���<�5��@���T�O@�Qr��H��ŉM�i�A2�L����AH;N(Z��?kҩ�v��"����A9v�	 ����E�Q�"���(�@#.�Z?�����a?��r���>�2u0��n@=p�j���b��C�9@��G�y@����}�A<K��ba��	�E�A,]Z@=|��[R?���T�����@ޢ{�@�#�PKH@6�N�=@��e��aA�ġ)����Wc�j��K�º� �,1DA$yGP,���ͩ�7]@)�����=V��?P�              @��X�M{�>�Q�q�c�@���	| f@��8�%wA��xt   @�8`uR�N@�x�bR�-@V|�����@y�dM�=�?,��?}Lڶ?�I:Z��@)�     ?��u�  B��d
F0>@Ǧ���A��,C�tݺ����^��"��A'`Jb�0�f���Q?���͒�a        =_<����?�2��%X�?.��is���a���üڼD��p���m��PG?T����)�=�A21�ΐ=}�!�؃�?���x�|@U�]��<]@�Ɵ�	>@y�dV�=�?8�ףl?�I:Z��?}Lڶ?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�%�/\n@�N�3�>�WS6���@�^����Y>�5Qܐa@��݌�-M                                                =�v�:��S@uvݩƮ?���4T�͡�uPhw>V��'0M?I��`���=�Yf��)?�̊�S�? D�wB_�}�F"5�=�k���9?	��Kª罪a�-V�q?�1�����5�т�e> ��`$g�>`��t�ȿ��ơV-                                                                                                                                                <�r��">'K�A䎣=��mC�I��#��-? <s^�=e�FT�Ip<�B����>Ah])Oш=�">�]��{�e��MR<m �I=��I|�I�<!|����&�F�!�4��>���~�+��(ݣ�G��S�С�>ni2E+9D                                                                                                                                                �%mAc�Tt>ꐟ�u��OJ�$��Vn(^�����ؙ�>qƼ�Qt��%l�B��L>���A�{>F����o>�y.�YYG�$�V!��=�n��ə(�?���CO?>(�jҋL���l l^���e�$~��b!����>j�u
(8�?����?i>(�]L��> �/ė�J> fŬ�?��q|>%P$�	��@&\��  >0��T�  ���b'�H���һM�$�`��Duɾ҃��F��@ >�B.  >6>,��  ?U,��w�r?���fz���-?���֪�f�mD��                                                                                                                                                                                                                                                                                                �>���I  >@�7� � ��������������ؾ��zl7�����!��@ȅ!� >C�k��� ?U-�瘒?���$�|�-@]���f�k��Vd@U|���i��I�4��2�>���M	�@���L�3>���G>�he��@WԿ��ʾP�ɑ,b��e,� "?����X��A=@��)�?�J��XP�T#�>0���f=���|��A��@��P���zc�f*<�P'D�.��cE�{N>5�''7M�#��أ��?���2C���)����2�g��;� �g*!�5=F=n���Gg=i��?�~���Ծ��޳ѡ�����iA�v��{�>&˂@<�?U- ޒ�?���5c�n@s�٫r�>C����@[�a��C�=����QoF              @�~��p]>� Z� @���	| f@��8�%wA��xt   @�8`uR�N@��T{�M@V|�����@�.S��=�nc
w<?2%?��|���[�`    ?ċ	�L  B��hEB �@�
}�JU�+o3F���`���������;�^@�.��751?���?��        =_��}��?���A>+?/��A��н��g��h��<	�显��Gmu?T�ݪE@�=�J�-B
U=~z��?�{����@UB��~�@�U`F�Ql@�.S��=�n���IN?��|��?2%?�      @/��[W>�                                A�e��@  BL+��  BL��                           >��g�./@�" �X�>����6�,@� �A��>�y�}�T@�j36C                                                =����C�@
� R0?���>���j%�E>V�\\��?J{�~�=����0�?�Z\�^pN?#xHx"S�v}�?�f=�2�/��6?
{ق����]ցk#?��ȣ�!�5�/D�G>!NA���>`{!�_'��Y7�˙W                                                                                                                                                <S]`p�>&��a�0=����䪻�A˂te�<s(��T��=f��%<r�mٻ>A2r���=��?kp)黁����J<l�n�'�=����}�,<!�/�⻾Fe�Rf>����ϼ��&
������6�y(>n�-�.                                                                                                                                                �$��9Yܘ>V{x4��Uh���� ���/���}3��>qJ�M�X�$�<�;>�Ɛ
N>E��A��>��-�'�w�$0�X�D�=����6��>�sBI>)!�7��K���[1̖T��eA�HMC�~�گ��>i�J�*���>��'>)!� ���> 3����9>�2�x݊�>�ٴC�4>%�#r��@&\�  >0���9� ��#۠y&��%��x-��a��OX�ҤI���@ )��  >6�ܣ=� ?T�V~f��?������d�,Hz�=?�f1�xG��                                                                                                                                                                                                                                                                                                �=k	%  >@�[R	� ��-����E��)�����������+uhz��@Z�  >C�TR�� ?T�a��?��Ř����,Hʰ� t�f1��Ham@TĹg��/�I�a�5��>�D �ik�@�1i=��>�[6�^�>�6+��B�@VQ@�����Q�G9���d�U~�[w����w�<A<H�GN��?�ҶSR#U�I݅��>1ƙ��=��
a~�B/ۥiG��� 
�M<�TBnD����z4�>5�@ۑ�#�zoC(?��ơ�Hm����6g�f�0~��f���Z�k=d`Á��=f��H�Y?��JIBڂ����T��+n-���(=�>'p��E!?T�Z�a�?��g���@�B>��>Cu[��z@o�mz =�H�'ЪD              @�w�F*>�%�{��@���	| f@��8�%wA��xt   @�8`uR�N@���R���@V|�����@��T�v=��6�ذ?��o��?��$X3+H@o�    �ğ���  B�1��(��@�HNy���*�H[g�)��˾�/���'�R��+��vtk?���nĽ,        =_���P?����F�?0x��W]��_���q��۽�5Þ�����m?Tat+�=�Vh��="�'v�?�����F!@T�M�OD@��g%��@��U�y=��|ʶ{?��$X3+H?��o��?�      @/��[W>�                                A�e��@  BL+��  BL��                           >��[}n�@��#�dY>��~/h�&@��Y��>�zg�L�@�OJ�yr                                                =���:�@
l��[�?ް6�NM����Qp�>VN��j�?J�7�@t�=��[��\g?��C6�|?&^;=���$�"��=���?
��X�i����6=T�(?Ћ �"��5���i,>".6�/%j>`��;�2j���å�(                                                                                                                                                <���u,>&k)��Ǯ=�	������j/���<r��C{C	=f��jz<P;��q�>@ǽp�؜=��
������ t&<l��r��Q=�F�#�0�<"�FUs�7�E�/�"�>����b����@���~"8��>o�gu!                                                                                                                                                �#�1Lm�>%M�I�����*�@���p�'�3����5��>p�0_�%�#�%(�9�>$�-6>D�s:��g>��X�_^8�#f���> �����=�R�~�O>)g���>�ǉ���c���EY�R��~|��	`>ih/����=�J\��>)g����=�����>�d}!7�=��n��?>&����@&\�  >0�N!�� ���*6�cm����A�c�b�c�ޤq���>�P@�@ �g  >6ޛc�@ ?T��Ϧj?�٬=X�^�+-�iq�q�e{`ԡ�                                                                                                                                                                                                                                                                                                �;x�  >A?��� ���U�
����n`A�뾩��+��X5q37�>��n�� >D͸�  ?T������?�٬��6��+-�;p���e{�M~i@S�^����J%S&�&>��;V�n�@����d��>��nh���>�j�L�j�@U��7A�,�QA��Hοd��o�����m2�A;-�Ώ��?�JH��;t1��s>18ū� �=���k�D�B�4d�ž���s�}<�^�;����
�l�>5���9�3�#���Й?�٭����\�b8��f2J��f���~=fq���!=f�I�T��?�oeT�MU���=��2��X-�����:|%A >(Eו��5?T��`��?�٤/��@	7�e�s�>C�,�6�BR6*V/b=-w�B�              @�Ȗ�p�g+��;@���	| f@��8�%wA��xt   @�8`uR�NA](D��t@V|�����@w{d�mx��R�Dy�?�Ls��88@*�Q��BEq1`�L�~۲��D����%�D��OONlD�:�ͺ	�D��(b��Dp\��Q&�Ca6�)���?���3�@�        =7�W�aw�>�Û>�2�?L�&렡b�x���)��� 1%�p�mk�a��>�fh���>O(�&P�=�Ȼ�#�P?vV�2K�c��i�I����6�ID�@w{d�m޾�R�!�@*�Q��?�Ls��88?�      @/��[W>�                                A�e��@  BL+��  BL��                           �A��=���HF�Q�R�@C�c�J"NAfW#2i��@
��G:aA]��� �                                                ���yA�N���BI�h���T��������i����>��?��b
��>�xak�0R?� �Gh��qQc�����]�zx�O,�&)P��?�x^��[>f)�j��Y?����7m�2#���b>�Z�h.C>��-H�o���&k��R                                                                                                                                                ���8�t�ry@��� ��.����R^���d�֘9��8S=�v1'��X=�Ƅc�>0��e��G���4�䅼�oS�D����GƝ>�9$b5���a�9">��'�sԜ>��eCp�#t���4�t��<���>��Ge�S                                                                                                                                                @S{�~�������ѷ��?��)%�����=q�<�ӨA8�������m2п��������?�ˮ�r�Z���^��V������Y10��-������?6V�R����9}��>?㕡O`N�u���^�����*L�>|5�ŗ��&o�}h�K�2��<:?��{sx%�=�wL�?��Zɣy)@$��y�  >��cj�  ?Y�c8�jU�����0��]�zp�oR�P"���������H�<��A��` ?�����0@�M�w�\8�(5�B�����J�J                                                                                                                                                                                                                                                                                                ?�S��  ?	@��  ?Y�/�g�����Jtb'	���#	�u��I,;Kf���u���+��<�?�l�Xa@�M����S�(6&{�����-��@߿�ޫ��@m��>���� 2'���@�m�������ńZ ��w�`U�A�Xm3@=6 �b�0�6ۥm{������P)A8�[��g@�P��9p@�	�Ef?ԭ�!"�_�����E�8?�6���:�~5�ߍ��Q�c�����{^�뿗���Ҟ��!7n�w�@�����I���A݋׃�J'['1A@c\|��?Q�����@����@�S��r�d�54�_4���ÿn�O���9Ft�v�Ҷg����?���>Jk@Ƀ�-c�A�8J�h?�UTx��@d8<�P=�F���              @��>C2y>�|�;D�@���	| f@��8�%wA��xt   @�8`uR�N@��W�@��@V|�����@o��hn=�;VJ��$?	R �s~m?�U�b�q@d8    ?��*j�  B�-a(_@���w?<�)�sfϵ���_��
����P
V��)q;��OW?���"z��        =`L	d?�io�r�}?1 6����6+=��ɼ�9�-ZV���`G|���?T@���q�=�`.�b�=���M�t?��J����@TH��H�@��螋K_@o���s=�;�ɚ&�?�U�b�q?	R �s~m?�      @/��[W>�                                A�e��@  BL+��  BL��                           >����I��@ߒ�w)�
>�nA���@��:��{>�`V��[@���m7@                                                =�+q�>@@	��J1\5?ݻ���~�� E8�.>V�	f}?K���=�!ў�k?�mem~�?(�rC(T�S��«�=��dEů?7��=�����L�?�E;��:�5��p>"���m�>a_%��x��>O�a(�                                                                                                                                                <jH��>&T:U=�:�ջ�+�n<r���W�=f�����<4�Q��>@�E����=�%w��Q���5ݶ<lB�e�=���@�<"�{õ�K�E�_b�}>���W������?!ļ�RԯΡ>p�U�}                                                                                                                                                �#=4e�e�>B�HB�����|J���J5_1���6���>pS/����#<���Ĭ>BG�"�>C�̸oo>�6�K"�f�"����+>����r��<�4~W�\>)�i8ı��a|	�q޿�l�P���}��]�>hmÆq��<�,9�ݮ>)�Zela=��(�N>�T
����<�|�
�">&SY�XX�@&\*'  >0���@ ��Q��6PO��C���"�cj�b��� V�@�EJ  >7+ ��� ?T�����?���ģ��*T�i0�y�d�uu���                                                                                                                                                                                                                                                                                                �:9��� >A'}�  ��[�c`,��G V��ᾩW%S���}�ȵ7�=lT�u� >DF�l-` ?T������?���X9��*T��7��d�sʀ��@SQG���:�JF9W<�>�q�V�@�N�G�J>�b�.���>і	�s@T�u��3�QxA;�~�d���^S���ۋz~A:T�V͈S?����3|���, ��>1T�#�V�=���ń�C]79�g���W��<�R7���fl_S,�>6,�M�m�#��I���?���hʿ���֒�e��S��e��)r�=`�D_p�2=c+_�HX?��q�ó?��!�$����}�������O_�k>(�fz*X?T��m��b?�ϼM��,@	���%��>DW��'#@BG�}��/=����              @�O]��J������o@���	| f@��8�%wA��xt   @�8`uR�NA��#�@V|�����@��kV��P���G��?�yr�2�@0}�a~�G�x=Eh A�)G�ʧHE�/��D	s���D��59F�D	��׌��DutZLQ��C2D���i?���3��Q        ��18��>t��Uj<?L�D��b�h
���=��;&��eR�0�l>�[N��V�=��z�ߝ%���g�S�H?���sE��c
�÷���\�[���@��kV旾P�˽��%@0}�a~?�yr�2�?�      @/��[W>�                                A�e��@  BL+��  BL��                           ��^Y�Tu��L�֯��=@2����`�Ak���{�@2�ϖ��Aa��w�[                                                �Uk��8����MA��O��QT ��L�
����ꍾ�k!�m?��j_��>��|4XZ?�t�]л*�g&qh(�'�}$A��JԻdS?�5���=���Ǥ�?�~��%�0�e���k�Q-��?#)gy�}������                                                                                                                                                �r,p�Ay���髓��TJ�%�&|�/� ��R�'a	|=�Y
k�<��0/��
>0��zQ�C��6�ݼ�襄��=�&wk�>ٰ_3��\�Ǉ��*�'1�3>�
tDk��=B,�e�4��f��k�>�M����                                                                                                                                                @Efm54�g
� ��$xZ��n?��v6��ǥ����ݥ&��d�@7z��0X���&9��q�� N�0����Mئ@}�8�w�>����E���,GCajY>��p�d�����5�z?ٹ��>T�w��N�#DQU`��>_�%�>�$[����ˎ]��?�f��`�>
>M�?=�o��@#���A  >�&�w�H >�f�������3����f�g�n�S1���fX�
pD滚|��Rpn����e����@٨��?f�&ML��ɳ�6��Pߊ                                                                                                                                                                                                                                                                                                ?���   >���^�G�>�ƭ�o )���/M}���	�$�*�	�U���=��
q�����Q������f�dZ6@٨�i'�&M�Ay��6��H��@�R��@�?َ��\����[ �p~@���ɋ]b����T����`C�A��b�?�5���i@(z��O�5��h��y��A7	0̰�@f��Vp<u?��
��_�?P�٘�㔾�w���[m?�lQTµ��&���7v�f���?ü�����#]���>���J�e�Hڴ�@�3�%Z��k�$,��`�;A?�@Za���r?����?��+m�@���ŷ��#�xRcZ�W�k#Ӯ��T+=.����g)YM��?+�]�@ʳ��ӡ\A
��Jw;@�_� P�@]�0>j��=�~��QO6              @��E��>����?@���	| f@��8�%wA��xt   @�8`uR�N@��.��@V|�����@�r�½=��'c�<?
	$��?�"������]�0    �����  B�pU�@����(�)k�����떒����JĶq��' <� l�?������        =`;`e�!4?��[ptݧ?1�nk�v��\(�L��ء�e\�0�L�?T���x�=�l�!�x=�#�5���?��L�@S�(&@�5!*��@�r�X�=��Z{��?�"�����?
	$��?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�}�0[�@�<����>�E�ߝ�@�j\��(>��^�@�a=X���                                                =�ת֏e�@	|
L��?ܣ! ��ɽ�W��Q�>U܉}�o�?K��&w��=�қ,<9E?��EՇ�?+��ivi��}�l�=���n?�,�8��k����{?�����D�5�lo�>#�h���>a�E(/������)                                                                                                                                                <�0FˣB>%��<2=�Kλ�(��K9z�<r�)SjN=gh����<��Ro�>@5($NH=����j��IPlj�&<k��^z�=��V>�S�<#��1B��E$���q>�����i��My���W�ײ~���>pd[����                                                                                                                                                �"�yUE�n>h�T�}���F2��{������9���MY?c>o��9�`G�"�"��>g`(u�C>B�*S�!>�~�4،�"�_20>`,�\ɤ�;��SO>)�[/�8F��2����̿�vP���T�|���}`>g�]�y��;��8��M>)�K���u=�0a��>>�3wGS�;�Emrc>&�Z����@&\�t  >1�@ �����w���l^Roƾd�>\Ծ���Pgz�`@��ܞ  >7��}�  ?TX�.X�f?��y��Ջ�)Z�#�bE�dO��3p                                                                                                                                                                                                                                                                                                �8��8  >AR$��� ��Ɔ��-��ү������=67R�Ҭv���<}�o� >D���5� ?TX��Sn?��z`bR��)[���R�dO�;���@R��]���J���^��>���g@��,a-�>��R�ݡ�>�˽�R#@T8^a����Q�]pv{�dX��r���ɑZN
A9[9�[]?~�CO@"�@"�o�>1x�� =�$5��3ξDP꾨��D��<����Zz�@k���>6q�
�bh�$	:�&/V?��{u�b����ȵX�e�,/~�eܓ��Y=g�r��A�=m$���"?������V���U�Qfc�Ҭnw�������M>)�@��s+?TX�3�R?��p���n@

�=�|%>D��.�ZB&�/�-�C<ڶ#!w9              @�rQ��O>���R@���	| f@��8�%wA��xt   @�8`uR�NA
k�3C�@V|�����@fR5��>Z$䏦��?�Y�G�NR@4�a;��&(��� B �EE�c E���C�C�Y����jĠ.ʻ��.��>K8O�D|4�)$�C@܈���?���3���        �"�<h+��>g�j;�Ek?L�V$��k����=�O@7|H�^1�3�=�>���J��>%-�팽�M��~�
? �<$��\����?�k]@�z@fR5��>Z$�F�@4�a;�?�Y�G�NR?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?��J���Q��e�@CkV,p$_Ao䢤�Ľ@C��,(0Ad�~��                                                >�:q$� A��)���?��O)/>A�.��Ⱦ����x�?�'�M8s�>���<�k?��o�U�a�`W�W31þ&?bQ7>�$�����?��/$��˽� �&6Y�?��E'myw�-QX�\L;���;���#?0���.�u�-#f�C                                                                                                                                                <�)q��B��	Я>��=���#aF�<]������ѯպJ%l=�@��ё=N����>/ؙ�w�;��:�+�t���h��lH= U]�uD>X��V<e6�G�B�&'s��[>�n�3b��=^B(�����,>�q�X�Yt                                                                                                                                                @��k�h�>�41|,��>X�hY�5��<E�*�۾��bs���%"&[@W�z�N>���4�/���c0�ܿ�y��m�@�i����T���n��*�fbMpx? 5�]L䌾��W���?����P%��5�u��?��N���>�aw�{>��'�Jnw>��N��?���%G��>[��M'߿A���&ϥ@"�QA  >����.0 �޳c��y��-$�Z	�p0wT���VJ���u�՚c̿��̩#���wSQ];@��j����$,Ǌ����C����O@                                                                                                                                                                                                                                                                                                ?�U���  ?Ӗ������.&�����Ci<�:!��TdR�� ��v;�C�̿��r"�[��wR-t��@��j�%9`�$,�I9�<�C��%��@�����?��]�^ ��1���	"�@�e{�����y���è�`�A!�훟3?��jՐ@|R�)�����dA52����@TjA1���?�7��-͇?W�,�� ��� <�g�?x��)�`��]-"4r:�9E���Y`��ӷ�wV`���R��A�M��*@�h~�JԌ��F!1X'���������@S*��j�>��p�>ٔ~��xz@����ٹ�tN��]�H�,�{Ғ�(��x�
���/���ޣ�v8@�����A������@1�c�y��A��~Ֆ=>2W�              @�q�!�������@���	| f@��8�%wA��xt   @�8`uR�N@����*@V|�����@fZ�6��9������?{�1��@�1�ۘA�IKB�� A�{>�� �Dw�۸��/��?'���yöC�N�C[�������g'`�¢s&ej?���3�X�        =mV��z>���au�?L��ƃ'q=%��r���ס�	���{.�R�ˈ>�$֗�{'��W��?\q=��֕>�(?k�+��?����e�?�rM�yU�@fZ�8־9�6t�F@�1�ۘ?{�1��?�      @/��[W>�                                A�e��@  BL+��  BL��                           ��&�/�"��a��R��Ῠzm�'wAk��!�s��f]B��AR�Wo��                                                �i�֗>��bI9��䐭x��j>%�+t} ���q��/:?ȱ���"���o �?�\EP]�?c������=��(�Ԡ�>ih׼��?)���Oԣ=�(uu��k?��(�Kx��3�[/zQ>��a��Ӿ��D�G����x�Ұ                                                                                                                                                ���H�qF�7j���|�r��}��<A�5m6���%�/T�=��^���y�Ҫ"Mr>BlT�=�s�˕gk<(g�`
a�<��Px5��=���8f?�H0�����)�ۍN>�m8�j�&25,
�=5�Y��>�H��raU                                                                                                                                                @3�V����|Ϭ-m>1Y�,"�?�V���6��%@-;��#��@�\*�0�s
�徺N�KK`�?����]W@���>��Zb����>���爾~S,��0>'�A�k0��fe	��D�f��$�`>�����k�<����wU�fJ\>s,�a?�lF��m�<	�׍��{��/42@%�;  >�c�S� >ĭ��=]���,�����Fyn����Cu�������p��P?e�䟢��?���d�W�@�np^�I�'�is�?�;ב�A                                                                                                                                                                                                                                                                                                ?���  >�1�V` >ļ#w����)���F����n�CˬP������#0?e�߳Cv?���ψ�@�nv�ƾ��'ʗd���?�>XEC9@��hڋ�g���h��쪾��P� ��@��XO�j��Gc#�m�!�3�,s<@�I�m^��������� �����ٔ�@맣A7���ML������?���q�3�>���Q)��a�jgZ��?^������1m�ݾ��r`��r�kڐq#Ֆ?lr�/�r�?��s���c@��Bo�.��mq�n@G=C`x�:-�5xm��%7=���u�T%G�@@rĮ5_�?ǫzv���BD�odM������N�?t�͊餋?;>@W�@��r��Ŀ@�/���׿���p�@A鐌�vi=Sla ޝ�              @�rn�6g>�#���@���	| f@��8�%wA��xt   @�8`uR�N@�/d�܋�@V|�����@f��:>Dq�z�;?r��6��&@!q��Y�ڗ�� A�ռX�kDX��x8�B��A4}�`���h^C"(k�Ĝ�D	�ʡ��B�'��K��?���3��        = �2���>������+?L��ۼEǽ?������{
�ȩ��}���?��H�:=��_���e=�(FM�ݤ?&�z�R�Y��P��z?��8V��@f�� �>Dr���9a@!q��Y?r��6��&?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?��;���T؇�M+&���A|ƸAan��4�^?�f�E�̎AI�1�,                                                >��~���w���%j�K���q�ˆ�����Sv����	�_?��s�u��OعPȋ�?�֢�?`2ܖp=ݧ11Z��>_�zd�?'Ex��ӽݘ�~&ђ?��E!�s1�4�N��ɼ>�]4��x�>�a8�(�_��>                                                                                                                                                <Ǌ�W�S��4<1�zU��XվH���Fk4�ռ�D'~=ؓ�X�ȼį�#��>@���Z=�
O{��X<SB��TӜ<Ԫ`B���=�;����B<S��JY ��*EV���>�-`'������qT�:����>��-Q=�                                                                                                                                                @1׿lQ�>ê'�$)���p6h�@ỵ���s�0f�+���J��
�ת�5D>����>����m��EOc?����X�xUMɘ.����I�os�<s0�Wd�����,i>O�<�lJ�Ѱw+�B�P��=��>�_j�I���;R�$�z�����$�@�>e�9��>��M	��;R\ ��H>MG_��P@&L��  >���(� ���~n�����h�o6&�5AՅ�9�:�C'�����ׯ$Y'�?N�(��?��5��d@�;��G���(+*��ږ?���b0X�                                                                                                                                                                                                                                                                                                ?�9��   >�Swt@ �ұ�q�9�������ԉfK����;Hݾ����������?N�XFnR(?���J�@�;�k�f��(+f��oH?���O�r8@�1�K2�?'7XqE^� ��Μ�@���-�`&�:�����4�ZVCj@��g5��fayo`����ʵ�K��HHL4�A8>l}���qD��?��񎑅^>��R���ܾ}��m���?q���"�ԗWۅ�p:,y��"�H���щ?Mh���M?r���@�^?�3����B����?�K �{�@>�����>��ܦ{�>��L׻@a�u��晿� %�:���;��u���1]a��?^4�ߌ�?�{���2/@��H�@��V�-��f3pټ�/@a�����=�Eh9s|              @�y��=�>���(�@���	| f@��8�%wA��xt   @�8`uR�N@�<����@V|�����@p����=��8`�!�?
�E^1^?���$���a��    ?�j&��  B�-�W@�O�38�(c�JJ�H���9�������DQM��$�;@��A?���}��`        =`_ >S@�?�-a�+(w?2^��������e
ӷ1��i�����P�h�?S�X�t=�x=��5=�u�:?��	H@S5:��@�ڰvdh�@p����`=���i�[?���$��?
�E^1^?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�!���@���e��>�&�&+�@�3�<l�{>����@��S�;�                                                =���r�@	 �y5?ۜ�hKƽΕ��K�>U�!Y:z?L!�(,x=��f���?�k�R?.e���IL�MB[�'�=�U�!�[�? @5RE��Ki��?�I5H��y�5�D�e>$ˎ]]>bd�SC¿�6�	?��                                                                                                                                                <6YD�|�>%6V&b1=�m��Ǫ���C-!t@<r]'X�	�=g��IР<�� �>?�a`�=�����d����h<k�KR�U;=�Eԛ�<$8y����D���Ra�>����$�ͼ�� �0j��a3��I�>p�hU��                                                                                                                                                �!��5�>�>����7��^8��S����`Uf��d'$�>n��E��!ӛAH��>�;���>A�D��I�>�ש}�w�!r�	o�>2t�V���:�)�m�>*<^��ٽ�
:����(�S���|q�H<,�>gW��-�:�4�q5>*<�vʛ=��@�Pd>��'���:�wc/��>'�:Nm@&\e	  >1;aU_  ���������`�Մ<��e�ܪ�ʾ�Hp�^�@t!�2  >7�!  ?T)02�	?�Ʉh~��(p��LW�c��|�j                                                                                                                                                                                                                                                                                                �7t �*� >A~��` ���]m$����c��%�'��Mn��18��ܦ@u���:��j"  >Dڰ�m� ?T)����?�Ʉ��l��(p���Կc�~.@Q�F�Fw��JƤ�"_>���f��;@�i�P�B>�^�an=p>�:k�� @S��w��G�RYZ���d(�dWɿ�ɜ���A8p�@��M?}�q�4H�b��M��>1�T�Q=��;�'��D�X���۾�Mn�	�<������(\"�A�>6����v�$2��m�?�Ɇ
�{��^j�̟�dx�'���d���&�=d#_!ʌ�=kG{�3�?�dA���r��O�����ܞir�`��/"i>*�&���J?T)c�g-?��zٹP�@
�����>EkZD_`BC���亊<�p
	+�q              @����fӿ�7��F��@���	| f@��8�%wA��xt   @�8`uR�NA�\_P�@V|�����@���%��D��ȴ_�?�"y���Q@7����w�A�4d�8B1A�)z�EJb��)gD��0�D����c�D�~GeHmDx8%蔖�:y�W�-?���3�5�        =u�B�~�G>`e�D��?L�]i�½�)��`=r�"���We�͏z�>�잧��>|Y���,�w�=�>�/����K���}��G	Bdm�@���%s�D��Ȳ��@7����w?�"y���Q?�      @/��[W>�                                A�e��@  BL+��  BL��                           A;8��]�kF�����;8d*D5Azt�=o<@br|��DAf���%S                                                ?�n��Ra�a�/V��?�&ݴ|L?��e�������W�@��z�-��tr��?��A�؎��T$c�.�?�g�V�1��,*�?�2�CЕ�>׽��G�)?����*(����]�,{*�ݢ?@_�@����j��                                                                                                                                                =�P�k�A�(z����=⿖n��=����)x�"�W� �3>*c.%1����4?�U>7Tm�$�M��*���ӌ=�a����b����B%`>1���Oy)W����%M�aS�x>�V��X�[=��6�����pB%r>��yL��O                                                                                                                                                @#���<?�� : !?����C����<U�Z�%�	t�s�����K�@HlJD�@��`V%�?�*J�@��aU���@L��`�fz@E��b�'�3G�R+�����7;?�B\�?ŢV)�C�G��@2���h��<%�@l�_�ǿ��4aX8)�2c�nR-?����|��@}ˮ�&��M�qX�@!�2�q  >��L�   ?��O��� ��!�a/�s�"�`=�W��ܴ����P~P��N)�8 A��'�|U��|@���,���"i�n�`���ۑ                                                                                                                                                                                                                                                                                                ?�n\@  ?����� ?�~�{b{���"�㨃�.�_e\t��#�Zs����~�J�bt�-T�&�N��G@�s9%\��"iMbt���V��ɳ�@�"<]��@���}�@V{��(@���;!�����qe^�G���()��A$���*�@��Oh�\
@��l%����R\���A3�����@�פ�6c#?�X���@�@]�H�?��e�2s忷�-�ub���Z�j��:�����D00W��@A���@!N�'� �@�|a�w ��Z\���,@yZ�q3��@F�B����
W��A,��`��N2j@��@��n@0�[`�M�@,,�Χ:��4�:l�Qv�]�����7b�@���P�fAģ&5��@CK��>>�B
64�zA�<��:e�z              @����6ᑿ�@�Fǡ�@���	| f@��8�%wA��xt   @�8`uR�NAtK$��Y@V|�����@��4��O�~�v��V?����P�@+�$�Bb���3��}� B	�y���D��~�D��A.�D���3)��D�H	���	�c���@�������$�P?���3��        =cS�Ye >�iT��"k?L�.t��������="\��f��kR���>����S">?��XZ�r�Č4Ք��?�g__?o]g`ӿЪ�+N@��4��K�~�v���@+�$�Bb�?����P�?�      @/��[W>�                                A�e��@  BL+��  BL��                           @ӎ!����z����� �ӌuB��A������@���>'A_(	2�                                                ?���r��'Ă{�ߨ?Ӊ�U�X?3Y0���@��r�)� @DjT�_��&� 0�?ԃ���R?kϡǈV�>�ۣߋÆ���+�]�0?o�k�q�>����L]�?���rNi��1�-�����;��?
��ֱ�I���خ�[                                                                                                                                                =���bF��D*)�v�$=�h�;�=PjV���-��"�+l��>0X�����F���Q�>J�ou��=���s��=M��_]4�32�=���=���A��u≫7�(���Ø>��)��D�<�|4�/� ����Ǜ��>�V����I                                                                                                                                                @@������?��A_�]2?K�x�1���j�t5/�+%ֺ��*��DfU�@L_�&��w?�4����?�$�	F,���o��=t@Q�g:H��?�����_�F�kp_B��m��E�?H���x���ݠR3�6�� _�x5�/������?N�'-�4�j�xCe$�����H���?�Ao�n�k�?Pt'ݿk$:%�v@$��WA  >��ȼ�  ?���+(���fU�2��`����VQ�Pm�����᎟������w�p��]�&啀@�@��V}�%�R��1�%T�����                                                                                                                                                                                                                                                                                                ?���  ?B6|��� ?���x�q��h�\����,(�����"N��&E��v�0�����`�\����ZV�@�@h����%��g����!��ͳ@ȴ�C�CD@gn(�>�@3�6}�@�k9R���j��n�����>��^A�����@v��	���@R��|e1v�����IA6nAd��r@�x��@]T�9��?���� �<?�����m�Ρ-��x �8�o̢�.���o#2������(�?�e!9M唿���0�`�@����Ly8��R�oG��9�Kp����X
>�t���2����c��\QO�@�My���u@1���?ݘ������iK�ie���1a���;k��@�П�/��A�h��`|?��Ʌ[��A�e�л�= ,�(              @���P��v��e�@��@���	| f@��8�%wA��xt   @�8`uR�N@�d�$��@V|�����@�æҙ�� |Ho�?f,�']��@Я�pl�A�d[�  A �����DH��?B�N��LV�5Zg%�Ccw=l;TD#!K�Ba�Tk��*?���3��&        =.?Lvf�>ǟՁ?�m?L��I�5��V�K�-��P�19 ���g��D�?XBa)�=����a=������?3�m������ʛ��?�g9� �@�æҚe� |2�y�@Я�pl�?f,�']��?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?���힁��E`�Z�ſ[�}4>��AS Y�Y1@?��w:�JA>^�����                                                >|g^^�.�$�.����)�8l�l`y���$��0�;i�?��~2�s���\�.��?Ȗ����%?\�7g0��=e�n��r>QU��Ux?%�l��}=��bm}D?�T�i�=<�4Ԯx��>�O���>ârW�H�7��(�                                                                                                                                                <�� �]]�1��F�{�,��H�#��BLY����݃�՜�=�l��t�R�2�w0J��>?�BF�=ұ{I��;�R��Mt8<ƅmV ��=����&/��/��'/;�*�/�
�>��9���N�U>��:D]N��>�y�����                                                                                                                                                @-�5��ft>���a?�������@'��|R<�ߺ�,��ى�'�mb�����%�>xы���'���z/�X�?��p3f1��_�>�G��#��:hRj��K��幩�=��j����#�_��31��>�"y�q�:����J�5�`��>U˞qyh�>��1E�,��:	&'��`��@@&C5�e  >��`�6� >����K�����{G�������/T|j����~S����?%Y�)*�"?��n��@������'���_�d��I4���                                                                                                                                                                                                                                                                                                ?╵��  >��+��b >���VhY ����n�ƿ���t�H�/�Rspc������A��?%\���<�?�a��z�@� �>P���'���sc��H˂��@��ۨΰ�?)i��<�~�"��@��/�+J��i��t,�b��@��x@�K�l�<tP�3$ȿ�NW��D���N�5�#A7���2�?�@2��?�6X���*>�:�X�
澲��Aގ?�n>{.�Q��1S0��!���߳����V�?&Qt?ӿ$s,,���@�(?�z����]K�.
���#�nR�@`�x�B>�/���ܾ�8�@Z$�{�F���[�Կ3�a�t��U�H��?5(��2?�x��
��@����@���ChjC?TCN�'��@SD  2��=������              @��7)ڴb>��?�]@���	| f@��8�%wA��xt   @�8`uR�N@�biu��-@V|�����@�8�m�=���=5�?\)m���?���!@SD     ?f��   B�[�v��@��)Fԯ�'�N,�4��A'jS���1n�@(��#Fbq��7?���A�%        =`nŊO�?h�:�r}?2��������E��$��Җ�s<��	\�!?S�2O!�=��,��M=�����?�?.V_��@R��U�[j@�^m����@�8��=��h���?���!?\)m���?�      @/��[W>�                                A�e��@  BL+��  BL��                           >эΡ���@޳g!�>����s@�
�B�J�>�R�M{��@��r:Ս                                                =��>e�2@��mk�?�Ե
��3���{M�u>U{�{VUd?L��X"�==���Ѐ�?�%U��Lq?07�#�{� �oz�=�/�ʶs?����9��y��<�?�ϲ��O��5�P̈́�>%���p]Z>bЬ��3���<Fw/�                                                                                                                                                <�81R>$�J>$=��{�#�����n=<r:3F��=h<*����< Q���>?^Yw1��=�㱚8��z��v<k���r��=��	�Co	<$��E��Dl!Z%BH>�����f���;O�����/�\�>p�H� v                                                                                                                                                �!O
���>�U�_L?��><r�#Y���R�fe��Yt9"�>n#�YeH�!N�L:��>��ץ7&>AR�x�z�>�[e>�t�� �)M�X#>�q��v�9��B��>*z������A�|����F �p�|c`n��>f���ñ��9��hՙ�>*z�0�=��'��KO>/�g����9�Z�F�`>'k^N���@&\�  >1]_  ��7�[Y�J��
���0߾f�w�B���nk��@@Ӧ  >8J7�� ?T���#�?��!�֠/�'�:���B�cJ��6                                                                                                                                                                                                                                                                                                �6nc�  >A�r5�@ ��A!-�������Φ����QpF����X��9�9	� >E�3̀ ?T���~t?��"[4��'�}ڀ�l�cJ��}�&@Qf���J���@R�>�VƈH�@�[���>��S8�>�.�萟6@S�s<���RCq��(�d��������:��A7��c�o�?}O��oپ�l�4�>1��-�{�=�(�k?9"�EZդ~\���:f�/<��l�2義����*�>6�H��엾$Y��B�@?��#y�8��!�ڛ�#�d
	|�F�d\6�E�z=pU-1$g=ryg3�?��e���	TG淾���3�k��/�n�d>+��"Ü�?T��o?��͚B!@
�XI_>E���)B�{9�#l�<���t��0              @��\l����K}X��J@���	| f@��8�%wA��xt   @�8`uR�NA(˽��@V|�����@U\�{ʃ�(^��Uh;?�
7���@D0kǏUs���%B@buT�T�EE��dJ�
,�%Y�7�^Dr�E ������D�Dw'a�����M����?���3�g1        =w	��P�>4pn��B?L�k���=��>ƒd�x�*�]ھ8|.vY	>�NO"�f��V���3�9>�;+�?>�fM�op�>���9?�qEzX��@U\�{�K�(^��V�@D0kǏU?�
7���?�      @/��[W>�                                A�e��@  BL+��  BL��                           @��Ū��;A�������K����An���]����r=��Aj���/�                                                ?d�B�h�?���2�p���mr���?&Bz��?�`F�z?��p��ȸ���o�b?��ㆿ�A�J���� 
>a�2���?z�Cr�;?��O�*�>�3P,Z��?�R��&>��_��BՍ?W�M_z0K���?|t��㚧��                                                                                                                                                =���|�=��(��Lq���H�e=B�I� �+=�"��)�=� $��)L����Fx�> aK�!��9�Z+%<�g���=����O�[>+Na]�ei�)s�]�վ��_���>��hh6��ϩ_��^�=�䃪�̀>|�e��"                                                                                                                                                ����l���?|�砲?>0�O��?��9�~�����T��?� �f���%�����?�6���K��OG���:�la��-C�{GT?�X�3������$����gߛ�M>��ʿa��?���ѯ�&"��-�?�k�<R���?���F��{����Of-v�N����˚�CI �L�3@�`_�@)�  >�$��   ?�i2�@�����O�B�����B)6��[}���)�t@�@TMU1��j@l�n��>�@� PrP!�5�ؼ@�ި�M7�                                                                                                                                                                                                                                                                                                ?�I�`  �ih���@ ?��Y�6����*U��(E��YS�?�E@�;�*,ؗE@TS��T��@l�/���@� M�t�t�5�Th@���z���@Ȇ򔼰��c6����{J�JX�@���<���@�JCݬ��2��)��A+r�h��������~�����_�w��H�<AnA1~�Ƕ���i��R��ΞeT�@8C1��?yh��B/(?��oY#9B�41���O@$�ˏ(���%aED@�Z��cBF@����1G�@�?s]��V��!�V@ߥM�J@@O�6*>ѿT����	���"��A%@��8�/@*�_�eϮ�񅚃�ǣAW��F+��=�R}���s�=vJ"���¹�EA��:V�'������A@0D*�=7UoD�g�              @��w�2>�>�S�@���	| f@��8�%wA��xt   @�8`uR�N@��1�k��@V|�����@T=i\��=��r�E6?����?�tX�q�@     ?�n��  B� �P;5U@����� �'V��|8���������=����!��x��<?��ƙ
#        =`�?X�YB?~G��츃?3���Ьc��j�Njdo��d2��˾�Cxn��?S����=������i=�>� �?���y6@R<�II@����ſ�@T=i\��=��I�?�tX�q�?����?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�,��v@�pġ��6>��K_��@���� >����͗�@���kL'                                                =��p�(��@0M��M0?��K2sl��G���b>UMf��C?MU�*��=��+|~��?Ǻ�td?1gJH�5��"��X-�=��ȞR�?��)����9k�FS?�?��eV�5��z�
>&���`�>cY$M5�c��ղGO�                                                                                                                                                <	O���#�>$����7=��MPXYl��Y��rX<r�W���=h�?*�"k< ˓��_>>��i� �=���񑯆��G��;~<kNIK�]{=��$��H�<%.�����D�����>��������$�̼٦Rs��>qH�ߌT�                                                                                                                                                � �zB�>�bg	����lm����9c<J��ǭ_�'a>m^R</�� �'�[*�>ܦ66�_>@���G�>�7��]\� ^�P�C�>�
�����9�>G>*�Mc���,Qy�e��Q�r�X˾{�5��[>f	��Uz�9�J&��>*�<����=����(>f��s�/�9?CN<�>'Ϧ��aS@&\��  >1�ܖ�  ����{�����)|l�g�k��ľӝ����@�g��  >8���� ?S��K�]?��j�� A�&�x��r�bȦ����                                                                                                                                                                                                                                                                                                �5=��6  >Aҭ�?� ���-CNbL�����[�����a�Nl��7/+�ǳ�8�#4� >Ek�ސ` ?S���
�?��k1�j��&�MKIq�bȤ�K@P�4X�봾KCX�⟭>�
���>@��5��>ƞ7>�f>�f�����@R�[�>�R���{�޿c��_�߿�ل��H�A6��n��?|��w,�<�-�X>1���s�=�ɋ�D|x�F�5�n_���bW�<�Hky�l�����mk�>7G����W�$�M��Sj?��lVU�L����_,���c�eL���d �m���=\LqAv��=o�9�???�����&�����ǩо�7&����v��@�o>,��/"�D?S�����?��`	{��@tw~�>F}����@��%�y==]E�\               @�r��%�>���V�S�@���	| f@��8�%wA��xt   @�8`uR�N@�Ø*���@V|�����@��:��A=��,؜�8?�]iFV*?�'�*[��     ?�ʄp@  B��p�xV_@���(v���&�,��������BT��q���g���^#�O?��ʠ��        =`���8?}1�Z���?4N��$�L��2߼�������'�Ͼ��YG�?Ss�B�-	=���H�%k=�O��0L?��r�0@Q�����@���Cr�@��:���=��B'�zC?�'�*[?�]iFV*?�      @/��[W>�                                A�e��@  BL+��  BL��                           >��de�@�5	׵	u>�ɛ
�#@���}>�e5��@�QNWه�                                                =�8�@����?�x��Lv��W�ÿe�>U#ns�~�?M���I�=��[��?�UA}�?2��	;��$���6�=�����?�P~���p=�'�@?Ͷ�&����5�1ˎ>'�<$3�B>c�^��R����A��                                                                                                                                                <	� ��_!>$*rF��=�E�e7��M FQ�<q���^p=i!6��gR<!G��wԂ>>O�O%��=�W�񇱻�9L>|G<kz�!y=�<d��=<%ʞ�PY��C�ݹ�R>���k��O$ɼ��^�Y�S>q���F�                                                                                                                                                � #��f	�>���o���p�[�0���u�֩��}�
JԬ>l�V'Q�� #VädU>
��)�>?��?��>~�
"5�D��P�L?�>a���E��8<�Yk`�>+e�Žƭ�F��N���u���{;��v,*>e��'�AJ�8<��"k�>+S��l=���R�3�>��,%2x�8<C�P.>(4-��%�@&\  >1�"�� �����SC��C̏5�9�i=U;s���σ�=��@��k�  >9.�� ?S����?]?����̃��&+}��F�bO� �-�                                                                                                                                                                                                                                                                                                �4 d  >B]W� ���������Fu�K���yMQl��k-?��7�7�S��� >E���w  ?S��8k�8?���U��L�&+��rAZ�bO�H2Mx@P;��`��K�%r��>���^#@�K���}�>�B���:>Ҡ���t@Q��0���R��d�F(�c����FX����3��A6+�r��?{ٗ@��� �{�.�>2�7�ǧ=�dK=��F��_�WZ��y#B϶<��<�iо����*,>7��.=���$��(
?��ր�=�����c��z�c�y�-�=ed�e,�=w3�yL@?���>f��{w6���k$��Q���'�K�>-�Z�Ii?S���(a�?��ɈN"�@�q�"�>G!+X��@E{�z��=zal̸`�              @��(S�V�>�}f6؎@���	| f@��8�%wA��xt   @�8`uR�N@����`��@V|�����@I��>��> ��/g�?�[�7��?����rN@E{�    ?�m�l  B�x�(���@�(�<כK�&j�]��f����q����j���8��xq�?���^���        =`�>$O\�?|&<a�I?52S�뽪���t%���y#y�����>�a�?SFՎ��~=����'](=��3ˮ�?���	���@Q,���x@�1� �@t@I��>�> ���?����rN?�[�7��?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�~��@���
|:�>��V��Ä@����-�>�D>��i@����i�                                                =�U����@^h�*g?�F(z�;��Ϥ�V��0>T��H9��?N#��^�>=�^L]��%?���e;�?3�A�
��'J#��/:=���@�?!��Z�V���?�A�?�3�H۴B�5�R�=�>(�� E�>drj�l]���kb��                                                                                                                                                <
���W^>#Ӊ�V�a=��(]f�Ȼ�غ�X��<q�9B#�=i��u�1�<!�
���>=љ�q�@=�gŎ(d��A�/�B<j�/�s2�=���v��<&kl}�0��CZ�A���>��ڣv��[ �����<ʀv>q�;K\                                                                                                                                                �7���D�>;k ���ￄ��z��b�M ���;���2>k��93*�7Z8cY>:��M�X>>�J;i�>}�����ܐ�G>!a��¤�7tj@��>+t�XZ��Ɣvm��ʿɠ�<y�۾z� ?��>e��E{F�7tb�l0�>+tΤEA=��УRCR>��o5��7s���>(��ɪ�-@&\��  >1���  ��[Jg�	�����s���j����~�����.��@o�>  >9����  ?S��m3ε?�V�9��%t]�����a�Z:�Zg                                                                                                                                                                                                                                                                                                �3CFV  >B5�͢` ��d��K��������(��B.K���Ӡ�_m�}�6�_��  >FP   ?S��n��?�Wqj���%t��g�Z�a�XXp�e@Oi�I���K�`���i>�ygi ��@����a<>����K�>��=5���@Q}��u�S<�/��c��?ث��r����A5t�K�X�?{2a;E(� �^n7>2;[�Z��=��c���G����ٿ��B.Yb�S<�S�%���+Y#��>7��E�*�%qT�y?�X��/��kJjE\��b������cgEY�6�=iH�w�=wgd��?�P�
�!^��D��A��Ӡ���&���H{�`>/Ll?S��ۍ�?�J�B�e@��V9lS>G���ehB$�%����<�B���a              @�8ż��b���w�@���	| f@��8�%wA��xt   @�8`uR�N@�kף.��@V|�����@����'�?�����G?�,��َ�@(В
���B"l�x���K��D�x�6���D�>�g��D����pTD��0K�`Db#:�Rn�C�q@,�.�?���3���        =���CRa�>�N�$���?L�������ן=�T�$ �oM��>�_��R>h򨤄j����j�� ?���W�X�2vpI�ĉYb��@����;�?������@(В
���?�,��َ�?�      @/��[W>�                                A�e��@  BL+��  BL��                           ��}��(]��0��qz�@���3QfAa�FC*�@G����q�A\��1��                                                �bȘb�iϿ�0����)Y³��Lze�b¿ ^��p?����l��?�F��I?����/�*�q�ƓNؗ��8s3�ȿ��|��?����g�>Ր��CZs?�S�"���2^&''����cX&��?2+LDf1�����^%                                                                                                                                                ��S��~H��B�����lV��y��!8�E����H��ܐn=�0���G=��Rކ�>0��.z���gj��߽DG�o��� �gӀ�>u�e�L�E ���*�;r�>>�Y]X�u=Y-ȿ����K^�>�6dFp�V                                                                                                                                                ?�@���D̿xN�O�� (�_��?�>וT�
�����fB�X�t�����	�ῂKKս�>�Ql�nAӿb�Bޅ5���8��k���du�>��(΋�(�}?�'����B���?��f���T:���M>�M�7Α2���d�j��@ܿ��R�\r?�Itl�ܼ�7�Y"w?����_@$��O  >�߭8   ?�엥�U���$���8�[R3m��K�K�Y���� �b�� �,������;D�.�@Ǚ5�\��#B(A՗j�To�Q��                                                                                                                                                                                                                                                                                                ?�4�c@  ?h{�� ?�՚ZDoU���a�$�� �X|��Pց��]��"n
G- �,��A���υ/�CU@ǙL�����#B_$53��T�^�Ub@�e|���@�#G�^�o�����@��j����Ě�ǧ>l��d�yG,�A�p����@�cg&�8����k����u�>��nA3��>��@ǀ����@"nR��@0r������-����?��ݘde@��㍊j'��$��#_OT���{+�4?�2{��_���̃&�@�:��>���~k�
��{�Wf@c���B�?����H��
��!#�@��\��C�.Ml��/, ��Z��e�	�1��8�.�p�.� �yW�>@�X�WZ/@�``c]>@=�}���@`�x)sZ�=��v�3�              @��0Q�>��>�~J@���	| f@��8�%wA��xt   @�8`uR�N@�+_w�FC@V|�����@��_!>�Qq�p?m�[V��?��8����`�x    ?����  B�^O>��@���*���&	�8��V��j�ޭ0��z��I�������k?����V'w        =`��N@�t?{$�~N)?5���lR�����T{ ��, �վ���FK�?S6���=��1��Q�=��r��$n?�7=lk0@P�\G��@��BDҨ@���)>�t7?��8���?m�[V��?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�1/��@��x���>�֧����@�nzE���>����Ͷ@��6�ޟ                                                =�@Q޶@��k�T�?׆\mJa�����~��[>T�vͺ�^?N�-��=�$�^8�?Ɨ'$��?4��g�ν)��)�~�=��줜�?�p���]�ug��?̶=^2��5�D8��>)��~F�>eM$�_��yB�Yb                                                                                                                                                <>\���>#��tG�z=��o[�6���vA�V�<q��;gD=j��7��<"G�RaS>=Y�%=���P��軠�YGaw<j�g����=�� �$<'�7��>�C�Xo��>��nd�߼�>v!+�����zc>r5�<�Qw                                                                                                                                                �8����>mː��p��0Epj���@L�=G"��6���>k`��w<Z�7�ls. >l���yQ>=q��ĔI>|���;l-�� ���>������6�>Qk �>+̔4��W���E�V��n���i�z� ��>>d�CP/��6�6�r�>+́�B��=�"R�</>qJ�ە�6��I$�.>)����@&\ TN  >2�  ��;!#�9����h��оl
.���x��7��^s�@#5��  >:*�i� ?S}��t�?����8�$�@g3�av�Wc�~                                                                                                                                                                                                                                                                                                �2U��� >BikSI� ��!�扡v����-H�_��l�)��ןX���5�iJ  >Fu��@ ?S}�4��
?�댌��$�z����av�k�v@Nj���L%QB�e�>�6�	*@����b/N>ŪZ�#�w>���c��@Q�#���S������c}�L�P�� ��E�A4�}.���?z��d��R���u^��>2h���n0=�r?z��L�H�%��Ô��l�Q�'<��j���侮d/-�n>8L����%Y�-�?��Ɛ~��<�=�R�b@$|caʿc(q���=n#����=x}�S�{;?�$�g���@�7��ז>�+T�*���(�>02��/<�?S}���$?��S@(�)��>H��ELBb_�<��H��              @�n��&੿"b��N��@���	| f@��8�%wA��xt   @�8`uR�NA)��@V|�����@3.�l�վ���K}G?�U���c_@0j�ۖ]B�"ӏ� A���GD���l�lD5�$�E/D����o�pD4K��ypDha�0Z�C"���0O?���3��7        <ّ�Q6rU>wrt+�?L�D�LT~�X�*�|��<��9�Q:<�el��M�>朾�a�=�r�˓���]��)��?����u�b�_}���%���@3.�l�㾉����-@0j�ۖ]?�U���c_?�      @/��[W>�                                A�e��@  BL+��  BL��                           ��>׬X��A@��@�$�_�8Ah<�����@GmqwAbk��                                                ��Y�������L�����.�'��P��؆���f��N�?����u>s7��>?��]C�ܿdF+����!"}
@H�݇��y2?����D��> ��5�P]?��\F��0�1�*�Ǿ��!2�?��onk�2�d��.                                                                                                                                                ��Q��opھ� �,���ÎNO{�6�lRE����
���=�����0�<���W�,6>0�ů�8Խ�V�.	Y��-^3�E�S.�P�#�>
�O�����T~O���*z6���>���x�s<��&88������nz>��ǳ�;#                                                                                                                                                @�~����7�e&t�gJ���X?���:�����_��ΰkyѿ������[��`�𾉵����.�n?�ྻm��oNM#� �Ѐ8����)s�kJE~>���Zκ���$��?��FЗ�6���V�MP����7���.|�a�%�����t���U?�҂ɻ�7���Z?]�:p+�@#�O��  >�{�|  ?��­����������fq�Mzy�QAbX,�՚��p��-�i��Y:�w�4@�����~�!��☬�����i�                                                                                                                                                                                                                                                                                                ?�x�p�  >ㄶ�n� ?w��{������D����[���_������a�ޜ��.�M7~��^��6@��ڽj1��!���R��xZ��@�1�?�p�@6EGU�ʿ��(zߡ@�S*
G#(���|F��g�$m0[��gA.i�ф�?����P�@�K�����V�SB8�A2B5Pd�@Y�0��k�@\���?�J*���~�,"D�aN?�9N�e�W�X��z,j����9|�1��W���=�Ŝ��1�y�����@�ʏ�0���A�}BO!�Q/�\d!�@X<�Tt�?�SFӾ���άU�@���a���'�0N��Ϳup!V%D��6�(���!�R����'`���@���$2�A'�P�K�@�Qɏk�@6t��k=l���BU�              @�r���B>�"�BY��@���	| f@��8�%wA��xt   @�8`uR�N@�aϐ$-L@V|�����@8����>,�?�?:\9a��?�ywݎ�6t�    �~���  B�d%��8e@�CZ�����%��� @I��TH�����Ꚇ������"W�?������        =`�>>��?z+}�n�M?6h���o����ˋ�FB��F�ܼ���pU�U2u?R����$=������=�6�:q�?�w���C@P ���=@�S����@8�����>'����?�ywݎ?:\9a��?�      @/��[W>�                                A�e��@  BL+��  BL��                           >��T��@ݦv��F>��}`O"Z@�R�i�b>�`��M�@��F���                                                =�s����L@��j2q�?��,��v��%�8>�>T�%�Ld�?O(��&��=�����$?�>��_��?5s�+g��,�&3��=�{]�?'S`�x���0�/\?�>zeF���5�	_\�>*�T��L�>e�c(hc���z�;                                                                                                                                                <�Xe��>#1�O���=�\�Sw�A��f��<q��SD=jo�<�`�<"�T�i=><�塬� =��ss����7��<j��#��b=�<|�,�<'�i�
���B���c�>��
�F����m �Zżܞ�K!�>r���ň�                                                                                                                                                �I	�8�%>�H�Zl��e��>��X�%H%���l?J��>j�9��G�Hm7_�>�t���><d#�ڏY>| ���Y����08>��J���6C��Ln>,'�5\Ͻ�n�j(?��Ss[ķ��zR��i��>d*�y���6<=t��>,'ҟ�=�Z�H�>>��f@��6�^�K>)jmxw�R@&\ �z  >2Aͫe� ���ke����9�Qv���m�d��о�nJed@�Gb  >:�ꮉ  ?Sd��@O�?�C�{v�d�$&_�3қ�a�HM&                                                                                                                                                                                                                                                                                                �1+u�q� >B��Y�` ����%�A��<=�͍ﾦ�M�y�9��(��q�4�R9t� >F�e��@ ?Sd�=��?�C��G�O�$&�2]u�a�S:4�@M{��ߙ`�Lv$�e�>��гɹ�@�@���'v>�k��,2>�R$�@P�,|�׾S�sw�hV�cdޛ\�ɿ�C�S 2A4&��(�?z�˫{+���O��>2�����=��*��r�Iv��K����M���}<�Z�ٸ�Ⱦ�����>8��%��V�%��ȿ9�?�C�/�a߿��^=�aᾜ��:�b� <U/�=f"m\ы=v��_� ?� WRz'
����������0�b���:�Ӷ$>0�i��?Sd���?�C�쳇�@��:Ʀ�>I@��c��B9P�<��C�%-              @�ß-4.���Ju���@���	| f@��8�%wA��xt   @�8`uR�NAs���6�@V|�����@���w�]�H]uJ{�?�;��my@4f�F�<B ZF� ��0PF��E Ʌ� �kD(��'|�D������D��?�(�Dp\Jd��C2V�����?���3���        ��]`
��>k7W�1w?L�U��cE�e�swG�=
�>�4��^p��_2�>��"�H*[=����LV�����i,?S��Q�_/�q�~g���wy�M�@���w�i�H]�)�b@4f�F�<?�;��my?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?�t>R��A�D<EB�Z@8vs~�}Al�Fl縜@8x�#�fpAe$pΨ.S                                                >)8��z",��]��E���	��<=�F��G����Z����?�p����'>�M��z�?����?�\���W<d�#����y��	�t�?��W�B�=ݘ�M�y?��E���-]ZT�S��٠g%SY?'>Nx�Q��
Ím                                                                                                                                                <Ef�f�$��
�|����c��<��_�)'��K*�%0=�	�Ae>a<��iG.��>0E�+W��հ@?h���H>dAĽ"5�Qk�{>����$�S�*l%�۾(��à�>�v�u�b�=P�_�(2����e�b�>�L�y                                                                                                                                                @ ���-B�>N���$��=���ɇz3?��"}VԿ��5C��m�?�������>dz�}l��n��e`"ɿt�F�zK;?Ⴘ�]�>�JKm6K�(�%D�>���;f쾓[��]?�L����� ̵'��o����8*��>��_a���SWB�H?�!���M�7�*��H�?6�ю@"�䟀  >���,4  >��WR�����I++ N�pg�'}��S�%�mo���π׊ڿ�8�v�@��．^=@דU�����;�� �8��"b@�                                                                                                                                                                                                                                                                                                ?��� �  >��sM܋�>ěA!x4h���H�@qd��⪩j��Ui4Ge:�����"��8���n���n�S�@דWͷՒ����$�
�8�q�8�V@��}�p��?�����p�o�~.	�@�un�k��X�-��]��ˡQ���AC&%�?�⪥5p@)�Ř�b��j1�?=�A0�X���@bxd]�T?�NX��z(?G/�ޭ���R扻��?�����	}��%���a�_o�Y�����*�Hg��pl�	=�@Ք�K�@�E�M@����i%m�J�Xx��Z@Q�هH�? -�ߣԾ�W���V�@��h8��M���z��Q�%�����n�2����`�P���T�p@�:屧�A4�-�@%��P�
f@>����}=t&��)�              @�ťeJ��>��7}Ӹ�@���	| f@��8�%wA��xt   @�8`uR�N@����j�@V|�����@�{=�>BґN?;��"X?�턁��A�>��    ���^��  B��HpU�@���0�%o�=�kH��I��v����vÚ���SG#?���h
y        =`����T�?y;�"�1]?7����?��H�Pbᐼ�����1����yÕ?R��*��=�͢ϔ�h=����z�V?����<�I@O9�OY*�@���
��	@�{=�e>B��"Bk?�턁��A?;��"X?�      @/��[W>�                                A�e��@  BL+��  BL��                           >լq�H�@݂h�%>��M��y@�9��Hd�>�r4�K�@��z��                                                =��C�f�@F��T-�?�(�HU���RbB���>T����e?O�:N)��=���V(<o?��ˊ��?6P����.��\�\�=�j���@?���Mӽ�Z쩨Z@?�����&��5Ϥ�>,�[�$�>f-������`���}�                                                                                                                                                <�;t��>"�/�M ^=���X]I+���g��<q�{�L��=j܏�p��<#Qy���^><wزk�=���ٵ8����E]"�<j��v{K=�����b<(U
�e!�Bl��X">����˼��b�����f����t>r�/Vp                                                                                                                                                �gͶ)>q>ض���'��B��M9)��D�������Рr-F>jH�����g2y�!>�ۉ���>;k��3��>{r�ʈ9���~$��>Ucq%*�5`��9>,���Vv��a�0����L��h��z_>��>c����*�5`����>,�℅��=�����;>k)B	���5`In(">)ՠ{/ܦ@&\!��  >2t6m� ���3�/ֱ����$t�o!���G�Ԧk��uB@��#�  >;>M�R� ?SO�D}v�?�mA��b�#��Cп`���@i�                                                                                                                                                                                                                                                                                                �0L��  >B�/[�  ���j���w���KK۞_���n�#KX��JJR_�6�4|v  >G;|� ?SO�q�v�?�mA�� �#�<6����`�����	@L��C��Lɔ��4{>����4��@��٠�>�5Ӹ��
>Ӑ)]O@P4�6r�T[\�֑�cO�����m`�	�A3�>�GQ#?y��8��̽�#��.D�>2�!PƘ�=�h�e���Ja�ڶ���n��<�18������>9)��0�&q�t5?�mC=��V����˱��a�^�d]�b��?�9=o[<Vmy�=~gxu��'?��23�F8����t�X���J@�6�d�nFp�B�>1���J��?SO�-S��?�m3#�k@k�A��>J	]���BS��6�X�=� �m=@              @�s��>��~���@���	| f@��8�%wA��xt   @�8`uR�NA �Vk�@V|�����@"'c�S�>X�*�P?���s�@9�Mu@���S�s��X�������E�P(��bC����,ĭw���ΔD���%��Dwp�r$wC1=k�DP�?���3���        ��x�"�5>\���i��?L�ad\��W�EW�Kq=
'�M~k�S�@ �[>��y�MG�=�>�� (��DƤvփ>�>���J�U�u�9�$?����	�@"'c�Sg>X��@9�Mu@��?���s�?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?�������E]���z.@9\�&sE�Ap9���@9�}G!�Ah#*�B��                                                >u+�=e�I���/��Ư?vl�<+>0�=�Յ˾�����c�?�bȯv��>����^�?��D�ڿUa&O� ��̕;��Ҿ�1g^�˭?����pw���$�&�?�Gj��`�(q�̑ľ߭[�r+?#�������	�gzݽo                                                                                                                                                <��=�����p�u
�%=����<L�1�Ԁ-�؄��φ�=�2�!�q�<����9_>-��մ���S���+����P�7�C���>�SQ�7�<b[~�*�)�&��v��>>��16���=T�N�ཚ�p �;>��#���-                                                                                                                                                ?��o�5�T>�^H&>E�;�Ɍ��*��=�<��kN{m�����Q�@���N>��{��p>\�L�}r����	3@f����d�Q+�n�%�����>� Rl��b6y�?č� �`�A���;��rɊS7K�8s�	�(>��(�ؾ��0�v?�C+�� e�8^��64��B��,�!@ ���  >�� C �҂٤����2���)��vOp�{�ݿV��Rv��F�O���ƅ�[F;��b, s�@݁3?���-�wP�4�e7(                                                                                                                                                                                                                                                                                                ?�̿   >��^� �� ��d�g��2K������I�Bq�V��MG�GG�ۙ�ƄΒ[�0��b,_MD@݁4{�-9�[z(�4�4��@�A�]"�t?�N�o6�@#��à@��Ё��rH���\����h>9A!��>bm���8�!�2GʽCK���6��H��A-ɞ����`�׌Z�B?� �hD�?(~��0ľ���դ/?K�W|������(�N���l����i�U?��O&��B@$s3�)�@�vC6^�����5@�|/@e������@J�_|����� <�T>��=�6�U@�����R�	)r_��ԿGE��n���MB��R��)�uT?�a�lB����!��1AꞂ)1�@)�Lƀ�EA�|i��=^,Ā>              @�+��F�m����g��@���	| f@��8�%wA��xt   @�8`uR�N@� �����@V|�����@=��#g�Z�:�H(�?x��rn�@yMFk��4��� ���L��JDUEjo_��CxA}�o��`����K~Ch
���C�JGf��B�?g~���?���3��        =��D��>��oG���?L�Xp1�m�45������}H�_<ܾ��Al�>���az�U=����x�{=��L�kI?!Yj�ٌf��0@	�?��.6ʬ@=��6�Z���L��@yMFk?x��rn�?�      @/��[W>�                                A�e��@  BL+��  BL��                           ��@0Y#/�QG����?��VI�G�Aaʀ��b�?��Xr�	AP�`�v��                                                �����&��VK{���Q�t\�d>ud���Aƾ��-/K�[?���cY�>R䴢��d?�O���F?Z�q׷�*Smp�-�>V������?$�h<=�Rη�?�e(���5�4'!�A4�>�D+�,�u>�7T������v                                                                                                                                                ��9�f6�-j�2a����DG�)<�&���D���?�E�eS=����S�S<ȋ��S�>>I!$��m=��)|�?���7�$<͞����v=�\o����iO�#Sﳾ-�C�L�>��(���'� �<����9x�Ṿ�>�Jئ�                                                                                                                                                @%�>�J_�������>��^lB��@��è��l�o�����yW���>���5n�����+J&������?���C/ �@T$�Y*���P��,��6U'���c>�|/+VC��/�y묿�ꌋ�e>�P���l>�ֻ.���5('�p���ax"HW���p�>�4P�L�5'�7�:F>��,���2@%�H  >�/��[� >��z�������)ue6��AŮB�fҿ>kݬI�e�����P� ?Q4�g�:x?��N�"@�0�}��8�"e���8?��Y�E                                                                                                                                                                                                                                                                                                ?�N];   >�J�i� >�g�s�˦���7Vs�Ο������>��F+����V�/�?Q0���3�?��3�wK@�0�H����"f%@f
�?��N��1@��1�ܲ�?��:��ſ��)ޡ�@�BZ�����0��f%t��,�h@🌽O��P��c�H����4f�R��HrJF�A2xYN��u��C��]^?�����P>�i��T������?Y�B�3ã�δy�܍8��F��D�Tu�m��?V����?�P�6��@�c�sFo���+�<��?��J�*3�@ �~mLl�?�0M�-���e����@jG���m��D��G�@Sڌ�@����]}Z�?`J��O?�H�x�z�@�߆�J�@�����Z��4|����@�P.�4=Q�����              @�G�Nxo>�q��-�@���	| f@��8�%wA��xt   @�8`uR�N@���7B`�@V|�����@ ���>rd�ᩗ?oK�?�c�W��D@�    ��S��   B��G��@�޾.��[�%4d'h���J��[�M��c�Lꙅ������Y?���۸V        =a��Wؕ?xT�9�A�?7�:
�����-'�����]���+i �?R�^U<�#=��k�=�ʢ~?���@N4�T�m�@�b�YGf�@ ���>r]��-�?�c�W��D?oK�?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�u�F�%@�c�,���>�7��X�@�%)A"�>�9-�K5w@�m�>]�                                                =�EE�U$u@��v
?*?Չe3����ЀӨ��>T�!8�~�?P�X��=����ia?Ř�=yV�?7 �~\�I�0�5.��=�Wp���?�2����܋�>6�?�^�:j+�5���T>-0���3Q>f�Z���=���%���b                                                                                                                                                <N5���>"�1�G�=�E����� Ɩ�F�<qr$�U�|=kG��I<#����><�C���=��b�q껥z.ݍP<jm!�<xu=�����g<) ��VʾB$���&>��֤zҼ�Y��t(��2I�*>sc���                                                                                                                                                ����X>P�����%x�I=��Z�	�a��~�x��>i�e��|
��L�I�>n�E>:���r$>z���k�����g>	֤T�^�4��?��?>,�8"�IԽ�X~ ����Y,�/��y�<��ɳ>cl�YA��4����9>,�#�`�,=���z�>���l�k�4�q/3>*AS�0a\@&\"v  >2�9�� ��d �j�:���Ү����p[����ξ����,�@+�KV  >;�yna  ?S=뛚u�?ٝ�O�r�"��*�{��`h8p��+                                                                                                                                                                                                                                                                                                �.�{��  >C��� ��m/�������������x�N(��Ԇ4�l��3]�Ng  >G���  ?S=�!,?ٝ��?��"��@����`h6hl:�@K�#�J�$�M��Z�>���ME��@����B�>��qRj>��6���@O��<���T��TmG�c=Ѝ|j׿��':��PA2�����?y=�|L��7��Ц>2�u���c=�߯�L��KV ���&���y2^��<��O�;<L��F�#�">9w
;�1�&f�����?ٝ	NC� �ߥ
�G��a9�pUNA�b�A��U�=l�D��:!=f�Q�Y$?���9U������X�@�Ԇ3%��]���>2T�+�9p?S=��o�?ٜ�?"Vi@�C�]>Jܲ\��EBwy�*�[=����[              @�m.9ؿM��b��m@���	| f@��8�%wA��xt   @�8`uR�NA���p�@V|�����@����8L������v�?�j��#T@A��&)��wr~���1�1f>�E'�gD���ć�,�FR���vZ�(D��#��/CD�� FhoQ�bX[~f�?���3��=        =1���3R�>FA#t���?L�ikY��=g.z����.��h㻾D&���~>��hg�*žx�MVR�=�Q�0DN�>�#����GՈ�&��?���+(p�@����7ξ����Snq@A��&)�?�j��#T?�      @/��[W>�                                A�e��@  BL+��  BL��                           @W�y ���H*̫�A��h���'/-ArR#3����Ze��\&Aj�خ�E�                                                >�yé7����\���?�4���V�>�^����L�6��Y�m?ѕ�u�){���!|S�?������M�DɣJ>'AY��D�?
$��K?�֟�p�>C2����1?�g�7W� 7a�,v�?�cZA�>�t]mv� �{�                                                                                                                                                =�����>� ��o�=�1�U�<�y�fܲ�R�7����=���g��"�����>)r���JĽ�w���9=<�6+@�#=���K��> ȟ�)���s�1�|�#LE�,w>�>�-�E���$Tv^�=��)���>{��h���                                                                                                                                                ?����?�k`�H>��z��/L�;��L���h��ǿK�<�@+�@��6x��?;�'�uUD?�K�0,����Sq^C�@!O3�W3�?���u�N�"�D��ȼ�]/�;|>�ؑ�8:�?�b�ؿ�2�`Z��[~?x���\U	�9��
�� ��c��y�>��?��?��ș���:�N�֜�?��	$�@"��  >�fR��  ?$K��`i��`'�g�n�~��M���W򈘭q��^YD,?�H�kM-@�P(�@�K�u�i��~�\f�@Q)�%��                                                                                                                                                                                                                                                                                                ?��>�`  ��jO� ?$i���F��_��5���'�!�z�?ns!�b�󡴯8�?���U�@����@�K��v�����0�\@Q+�����@Ǭ0-��'�Z�w?�Y{�l@�K����@�di1��F"H8���A$�c%[�1�3���p'^�Q�򬆧��:{�>ڴA)��-�n�~�
\�q�����v?���̆���o��X'���cP��"[��8D?��Mv������P�-@$\}�%G@<��4@�'g�Jk��D-k�a@l��h�l @B�-���\��t2en��2��}��s@��jC��@� ����<x`u
����E3iv�?�A�~��{����#Qo��?&	���AQ�hl�k�P���T�B&p����2=P
�O@)�              @�m/�a^ܾ�C�M��@���	| f@��8�%wA��xt   @�8`uR�N@�ب����@V|�����@���;M�@c��<�?���>1@'+uƒ�B%���� B=7�䱄D���A=����H ׅG�~K[,���C!⡽ǭ�>�lp)v����k�=?���3�fd        =`���-�>��4<@�6?L�X��=%��]F ��颸�Bp�q����>�HF��������+��}=�H��1�!?�����?��L61t?�ccC�@���C�@c�fL@'+uƒ�?���>1?�      @/��[W>�                                A�e��@  BL+��  BL��                           ��E$��
$�e�(�I�����(@(Ar^���Ň��b��%�A[$B��                                                �We��_J��C�q\����
�t�a=�No�m�O�ݏ?����?�Q\���ξ&!_����?��u�C�e?eM�R��=�N����>p� ⑄�?9��@�=֎���6?�ʨ���2�#%�3�>��1�p����H�j��H�֟�                                                                                                                                                �sٯ��ɾ6H�<���Y_ϛV!;��.>�4��"E���=�ߠ�������9�Y>B�:�n��=ۭ *(�<W�~���<�ǻ�n�=�I=$��M�Q���׾,�L�rS�>��#L2'�,���=C�t�!Ӆ>���g\�                                                                                                                                                @0>��*�X���0�j���0�}?Ԫh�^���IO<!M[��G�Y_@%�R�ɝ�`
���O�����%�h����[@&@i�~�عn��O�;W�>U����,)!]��>Q��
rw��,��6ݫ����s&v>ߡ*��;�5����]�pJ����.>w�%�'?U�[4�3�5���z뾁�Owfb@%�Y�  >�͡IAX >³h�xE�����?��G�XK�(�He�s��{��Ii/xߠ?x-�*�P?Ǘ'��@�c`tA�!1��fVX?��ji�O�                                                                                                                                                                                                                                                                                                ?ۏO��  >����A� >��}��c����Sס��[���H��'�����J�l�0?x-��#��?Ǘ�wf�@�c~ՕV�!1��+��?��d��@�HX�ޘ����dcо��ڶ&�@�#*�C�eB�R]�P?eu�����A���4�:����R7[��W��7�G��jʎ�A1dR�&��
�S5��?�e��쾰�uF���>2��e՚@�P����v��QeB��?2&�:����+���?|�}�ٟK?� o��@����Q���ƐV��<	?߶�MV�J�s�^i������}����J�Z�@�0���??�@�K�X-�D��݉ ���ge���?�E� �?��K�n�@�k��^%@�o7)t���A�A�!�,۷u= ��ᤌ<              @�mzu�����G�e!@���	| f@��8�%wA��xt   @�8`uR�N@�q��a�C@V|�����@���R_P�[W�+?p`T�7@SvFfil���O  A_,���DD@�s�	YB����,�B\�=s�B��;N8��DP�l�FBc[iCA��?���3���        =$f<[�n>�]��F?L��?P�N�Mp���K>��u���~=���� Xb?�zg��=���z_�=�ƹ�:�2?*����o��G�\I?�s��@���R^K�[IǦ@SvFfil?p`T�7?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?��¬��C����7���׋AV ��G.?���B�d�AF��M�F�                                                >�v��1����0�u��̑��HȾdiX������?F��e?��6M
%�=����i2h?���y�?WZ���=<��^�>T/y^�ѽ?#��
\��=�����ڽ?��m�1�4�,�6��>�՜���>���2a�d��W~��                                                                                                                                                <��ѫ��C�):Lz����HJ��Q=L��3���lG? =�Hs��X;��=а! ><�	��-�=���f¹;����'�f<�96�@f=���@M��&S�����.ep��">�VK�c���Q �{)7�@h�k>�U��C�                                                                                                                                                @"c�݌�>����,��y�!���@�x#W�¿�9h^�����l��>��}ߍ<>s{f���۾�	fB.��?�Ǵy���B�E�k�_��4�C�����6�:;�<=�tU�ݿ���q׿9�d�rE>��&�H_�4]l����5���͉w>T��q�>Ԓ�.x�"�4]�ਵ�Z,t8�݀@&& 6�  >�#���� >���s4�������04��4LF�����d;�� ?7���}��?�6�@@���z�"9�厙���D\���D                                                                                                                                                                                                                                                                                                ?�� ��  >���Ҫ >�e�������-����0Ɵ峿4ir��c]��o٢ؔ�?7��R�S ?�5�[�h@��r8vf�"9̭Aew��D]��t!@��9�7��?
N-GN�.��<��<�6@�zts�b�A	r>��9+��S4
@���2�P3�Q�
ڑY<��Th�?a,����  B�A2B+yȭ���qH�8?�.��sɇ>�~8F�28��Ҷ�"?��/�̶H��9Ǝ����pm=y/�/���]}�?8"qCf?16�#�{@��A�+h��\����3?�H��$�4@L�9d�&>��R�-�xYC~%g@Z^X�+z����|��5�v]`����*�`�x?G<TNQ��?��X0k�@���?���@�w�P�V?ZGF�O'�@�!@��i=F����JX              @�g�S�B>�Tm��@���	| f@��8�%wA��xt   @�8`uR�N@���æ�@V|�����@��kC�>���/Gj?ڑ2븈?��@"�I��     ���!�T  B��y4@��j����%d>�)1��V�'ғW���������;���?���r�ؐ        =aAՎO�?wvb���+?8��Z�vv���&<�E2��a�fI���#0b�?R\7����=��5�&7=����"?�_m�Z�@M3P�k@��
��@��kC��>���8uY?��@"�I?ڑ2븈?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�G��@�JX���>�7���zt@�l�aǅ>�	�����@�O ���o                                                =�ԇ�{@��a�T?��X HĽб���V$>T~,�"e?PRPG���=�f��5�?�Km���?7䍼�b�1Һ[$A,=�G[�'��?Qy8�w[��^(�E�a?���j_��5�i���>.d3��~�>gc��"ȝ��Bo_
�                                                                                                                                                <O�Xg�>"Yv>�=��Qf;y��T3Β<qb����f=k���%�H<$e���>;�^�]e=�
0�\��'�F�7�<jX>���=�3�m
�<)��ᚯ!�Aީ�8�->���Gӛ��$�p��n����%'#>sd��^(                                                                                                                                                ��f����>L�A�/Խ���eR ��+	�rS���`S+pr>iY�A��K������c>K�A_�>9�2�9�">zH����]���P>	(�5�40ـ�}>-E�:�Cz��R� l�6��v�	a?˾y����>c���^�4/��ҍ�>-E�<�\.=�[���>�8>���4/��E?v>*���`�9@&\"��  >2ݜ۽� ��0/�#����Q�n*�m�q4ZJ_���b�H`�@�Кp  ><m���@ ?S/^y�!B?����|?U�"wS�����`�I�%                                                                                                                                                                                                                                                                                                �-jy�  >CIޤ�  ��9Xm1����S���R��� �+I����}���K�2�y�v� >H·G  ?S/e3�?���N�=`�"w���<�`�7�,@J�����My+�X�>�Na��t�@�W�Q?��>���g�>���t�@N�TujV�U1�\���c/A�>D������7A2w����?x�=x�Xؽ�S�m��>3.����=�MdL'��LS�I�ƾ�� ��v�<���Ւ���`6���>9�U$��&��R+�?����0���u>�5�z�`� <�)o�b}�!=d�O��FS=~A�P/�<?���R������]Ǿ��s=h����� ,>3 2D�6?S/X���?��֡�Rh@�v���@>K�w��@N���L=�~!W	              @���*�a>�1-��j�@���	| f@��8�%wA��xt   @�8`uR�N@�ZG�{��@V|�����@ ��5�>9m��ó?^��[�^?�pQ�LN�@N��    ����P  B�q�T�W@����6��$أ�����tg�g���ۈO��\��w�T?���U4F        =a��2�?vtפyd?9_E�ɽ��j8���X�)D���ݓ��p?R!U����=�����=�i]��,D?��}0#D�@L�1(@�tq/��\@ ��6
�>9cy���?�pQ�LN�?^��[�^?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�O�M�@�2c#�4>���gw��@��ۘ�>���fN\@�1�q&�                                                =�8��`�$@C�PY��?�I�Hg����;3�>Tm3ث-?P�q՝�=�7�IL��?��m|�NK?8�1< ��3p8�
��=�8l앦?���+��� ���?�}[�4���5��o>/�}P꬀>h%*T��A����R                                                                                                                                                <��m*�>"
�#j�=�6Lx���E�<qT���Sb=l/���w <%t�P>;6{�ɐ=���&Xr��@�Ζj�<jD��K&�=��o
��Y<*�T�D���A��9i݉>��rw�R��!������P�>s���?M                                                                                                                                                ��X���>�/*(gý�����^���nt����C�xZ�>h������1tv�>�;E/! >8ɀf���>y�*�_���oc�+>
��W)� �3���7��>-���x&ؽ�P������zW�59D�y�It��>b��8�3��X�!>-���L�o=�@��[�>(�lk�p�3�A�L�">+7k#�@&\#\*  >3 j-I@ ��+�H��1������rF����g,��0�@`bP  >=3=�$� ?S"��"?�,�vB�!�5O ʿ_�����                                                                                                                                                                                                                                                                                                �+�n֎  >C�Cj� ��4�; ������e����+Iq<����#���1�P� >H��1` ?S"x�?�-7mu��!�g!!��_����v�@J�%׾M��X�\j>�I��Yh�@��)���>Ľ��z��>�_ַ��K@N3��$�0�U��+�w�c!�ԞLL��O}onA1�i�z��?x!�'���L!ķ��>3o�<�D�=���z�M��6�����+q�z<�|u3�4���9-� >:m��P��'Y�㖤�?�.�5�ڿ�I�%1 �`����qۿbah!�fq=gcsLy�*=��@>?���=Ͼ���Px"ھ����)X� XP���>4%�5l_u?S"Y1�!?�NH�x@W+���>Lا�I<�@F�P�S=0���v              @�1R���>�"��Q�@���	| f@��8�%wA��xt   @�8`uR�N@��36r4�@V|�����@ BoKp�>	��߉^�?Ι�Z$�?��V~�R�F�P    ?�7�Ǭ  B����/^�@��f�w���$��Bp������f��gB1m���Z<ή�?�����        =a'�e�J�?u�]+dD�?:��Y�k��B�e7������:���No��?Q���
Q�=�w#��n=��K�J�?���f��@K�\Hw�@��`����@ BoKQ>	��e�?��V~�R?Ι�Z$�?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�4E|i>@�#�"�>�Ⴒ�]@��L�+�%>��j��m�@�p3��                                                =�c�e�8@�oQe�?�Ŷ�.���%g%��>Tb�2�5?P��H���=��ve��g?Ĭ0 u� ?9n��4�:P;��=�/�Wә�?���8�����wj�?�>� �5��Fϗ>0������>hȿ���߿�3i%���                                                                                                                                                <�	�>!�Uy�o�=��i�<�t��1���<qK��G�=l�UߐU<%��y>��>:�;�@��=����)+��\���<j9r���=���B۱�<+3�g�z�AO�K�.>���:^����_����mnk��>t�Aj�                                                                                                                                                �;bz9�>�*6������1����8X.�辡2.����>h{S�B�:����>�-��Ru>82�+^B>yBel�Z�����+>X2-�v�3p�ي�>.)-�4���R���h�¸�I��y��3��>bu��_3�3i�橾>.)-���=�*���3>�?"����38
}>+�uh$�@&\#�  >3Y�35@ ���Wf�Xm�������s4�E�2��է?X�.@��ǀ  >=�϶� ?Sd;�v?�_Ǭ����!g%Dp�Կ_�                                                                                                                                                                                                                                                                                                �*Nn�  >C�[�  ��y�s�����F��#�����E��Q]E�V��1U�J� >I�Yˀ ?SjP�|?�_��)M�!gU�&���_���$@In�o3�NH�-��>�0�<U@��^|�>ħͩ��(>ԣ�.�c�@M��k����V6<��*˿cCBڿ�_����A1gX:�Y?w��}<ܽ�y�74�>3����=�5[r�O��N����٥����ߔ�9<�s�&�
����H�~.>:䘔�*��'��Դ�	?�_Ɍ�'��0��	��`^`2\#�bQ����=p �+��=�q��s�?���g����̩-)���QQ����� �����>5����?S\��ӗ?�_��DS@��;��>MҲHU��?�w�AL�<="�gu��              @�p�Z>�RH(���@���	| f@��8�%wA��xt   @�8`uR�N@��/���@V|�����@ �'�7�\>9��K�?Xp��-?���ֹp?�p     ?�{��  B���?��@��S�����$���>5����������0�0�A��?;@5�?���
�        =a(�O���?t��8���?:�Ŋ�	ν����Ge�����ƾ�t���9?Q�����b=��̩�=�j���?�:Tv�@I���N�@�j����@ �'�7��>9�:��?���ֹp?Xp��-?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�U���
@��P�@|>�z�u�j�@��K7�NM>�2�X�@����5�                                                =�7���I @���ї?�/�P�]��h�Y���>TZ���H?Q ��d�=�1����?�[+��-�?:1���"�6x-���=�)J���? �dm��-u0��R?ɰz����5�� 
�>1\�Ǔ>i����ֿ��fȡ�,                                                                                                                                                <M��B��>!����w�=�GM���û�j��-_<qE G"a=mo{�<&VS��� >:q�I��=�����0�dUn<j1/�Dz=�?o��$&<,�c��A)��>��C
����+|e����"
J>tZ	�2��                                                                                                                                                �t4y)�>'��J(���Ë#H���������$�5x�">h긙�Y�s�?�}N>&���>7S�h��>x���$����t�>6r����2ro!���>.���=@��Y�T:��������y{�5�΢>b(`|��*�2rh ���>.���Oo=�\T��>�46��R�2r@��>,5�����@&\$��  >3�U��� ����A���l��{��tb���ǫ���l%mRf@�4z�  >>���_@ ?S)ז{�?ں/��/� ����<�^vv�跇                                                                                                                                                                                                                                                                                                �(���  >D �?�� ��A#@!��nmc�0�����P�բ��G�0�1ـ >I��_�� ?S/��4=?ں��� ���$	ʿ^vr,v��@H�hW��]�N�o
�>�����@�q���1>ĖN�&y�>��`$��@L��f>C��V��(F��c� B����?+�#A0��i�Q�?wH"*�C����5�>�>3���J�=��G����Pc_@5�����2<�3�X�^��,b�T�>;|x�5��(xJc�W?ںz����%f���`�)�ֿbE�k/��=k*G"x:�=��F�9�?�C��D���;�\��բ�Ga��!7~�1��>65�lk�?S!Y� ?ں!mH@6]��>O���yB��_��<�̙�|��              @��f�I�������f�@���	| f@��8�%wA��xt   @�8`uR�NA �r-s_@V|�����@ ��6o�H�?t��j?���c*�@/��6����{�b��A�m|��D�߻J��D��P��jD���[ݐ�D����P�D\7�FC�������?���3���        =h>����>{��I�?L�A�ty���H-��鼷2:�:� �f>����>�	���A>0^�Q��=Y�8�� ?�{��5��_X�OEk$��f�n�H@ ��6o�C�?t��@/��6���?���c*�?�      @/��[W>�                                A�e��@  BL+��  BL��                           �{�B��p��%�$`K��@|3�z���Ae;��@�tPD�Aa�����                                                �)�Mt
9Ϳ��Rő���������Ոz{^	���9^P?��ƈU0>ح��P�?�e�gKx�b��1Eu�����0n��U�F+��?�kH^��>�"�;H!?���g���0� �C����wµ�K?���g���9��ծ                                                                                                                                                �F��P�����;�K����"���|��D�^e�~��ی�5WB=�u~�V�=PY�f",>0lSբ����T���褿��gG��G�> K�34�]�c˘�-%Y6�u>�H=r��=4� 9@ �|�j�]>��YW�Y�                                                                                                                                                ?�R+����=�p����X���?������@
��]����/���,��qz�MK��K�>��.����i���|��)a�-ɿMt$�T��&��s���?G��Vֲ�,���?Ў.E)����a��E�Ó��RT�3>�I�L�*�e B��r2Au�(�?�xl[�^�2�����?�0���/(@#�ٮ  >��㝀  ?���C����� �!��eo'׮[Y�N%ʮ�]�� @Q'�ֿ�n�Z�+追4�镺@�0p0t7A��)`���q�Ǟ W                                                                                                                                                                                                                                                                                                ?�J�   ?1��c� ?����_�e��}�X������,K׿ñ�[��0� Ax�!n��sf��Ϩ��W;����@�0y�60�ҁ�^���x�@؂�󐥢@�������F[�����@��k�W����ݯ��~�����X��GA�Q"mA@ft���U�\=ש�^X��r����
A-~�AZU@����~�5@&���?��K放�§��Is?�{[�����v����b�>��C�g�jI?�8;SYO����B�n@��%v�=��Q%;�}�7�-�CTc@V�@�&�r?�oeE��u�x���4@���;,��0��M�H��R���	+�0�|�����?��+?���n@���Nxp�A q��=�@��[��@ �.�N�=WO�
צ�              @��ewhC>�V.m�@���	| f@��8�%wA��xt   @�8`uR�N@�.p��PH@V|�����@ ��F'>�{Nvs�?�x��e?�	o]�Ε� �    ����V0  B�/<�#�2@�9���n�$�-vL���=����I,�
]S�#����?�����J        =a(�I��$?s�ݍ�g�?;���»���L޾W��!-�3U�� ��l�N?Q�->�A�=���f�h=�I�V
��?���wc�V@H��p݉@��"�x0�@ ��F&��>�Z�� ?�	o]�Ε?�x��e?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�N�1��@����:>�2�^���@��\�->��E�y@���J                                                =�a�3h�@c�1f�(?һ�;:غ�Ѣ�c��f>TW���<?Q[N�}��=���cz8?�g|�@�?:�#κ]�7�B�(bK=�'wpFB�?Zi=������R�cA�?�Z
C#8i�5ֺ;��>2O���g>j=�B�������                                                                                                                                                <���x�H>!LU4�W�=��rn_a���Rd���<qBn���=ms�{j <&�<�_��>:$'�+=�f'n8Z"���0�DY<j.�̂�G=��C�"|N<,ͥ�ކ�@ͻ֣�i>��Lzi\�����f��d�-Gv�>t�g'�	�                                                                                                                                                �ٺa��>lh�Sm���!�������#������VZ>g��]����#G��>kWK��>6����>xx�������2E�>�_�\��1��թ��>/5c�߽�c0a��j��:(���yx�|�/�>a�y+���1���nX�>/�s�8=�)ЈR(>IP��q�1�?e�s>,�,��>@&\%'  >3ކ@@@ ��p��[3w��/����ug��k�}��;זV@Qe�  >?{�.�� ?S�
�?��ڴ�� v���^	`�h{X                                                                                                                                                                                                                                                                                                �'����  >Dc]��� ��uI��'��1�<������S�����t�����00z-�� >J1�+W@ ?S�r��?��=��i� v�>]tۿ^	\��T@H��1��O&a�ֵ>��;�@�4�d��8>ď1����>�@���@Luj 2"�WV�do�c��5l���,D3A0v޻ �,?v�㏡槽���z��>4*A����=���.I�2�P�_�����������<����^��8�M�ݬ>< ��6�)� ��#?��֕����6V���_����h�bC� qXx=o��w��=��25/2s?�` #nTھ��z�3����g��]��!�bEtZM>7:��["?S1R�?���&�@�AA�a�>P�߁��BBc*I�=@���Ue              @��ǿY�9�@���	| f@��8�%wA��xt   @�8`uR�NA�6s�[a@V|�����@ �j��^�xr�i��?������q@4	��<*BBPE�뇐B
=!���D�WF{�ˢC�Y4^D�`���gRC���Pq��Db��2���C OtH���?���3���        ���%	�r>o�/�!�?L�U��Z%_}���<�>��!#�_P2�g�>���ZQ3C=�A
���-���Oc?�K�͛T�`H ن�ٿ� ���@ �j����xr�<ns@4	��<*?������q?�      @/��[W>�                                A�e��@  BL+��  BL��                           ����F�p��8����c�@'
>+jF�Ajx�N���@&KX3��Ae{v&Pi                                                ����������g����O��]T&HF��4HB�R���8�}� �?�RrM
��>wtk�؅�?��T��yA�X��E�uʾ�ð̎��s��K?�J�{$�>����?��멱�z�-�)bھ���b��-]?ؤ��\��	�F��X�                                                                                                                                                ���.3�~A��:���;���*�]�ȼQ5+ y��8�}�9)=��_�%�<�x�}ɢ>0�|]��0��i������5tx˽?�,e�ܕ>	�-�����g�+��MfV>��;@:=4kB�[�ݽ����D�>�3MB��                                                                                                                                                ?�3zyY����J����I9�׵R�?�@>Ӷ������-Yy���T*���� BLg���TV!����ۊ��A�iDI��� N��;���i-��&Ŭ�Z�|>�: �-��_�ٶr^?��Ȝ��;� �-Qc��5�k7;�|�3s�M�#I>��_Ȥ�������
�?��6����3/$����?I��o��@"�e�  >�Sh��@ >�������v�AX��o)P�Q��w�����5�����kK[����R��a@�����\��"-!v���%�����                                                                                                                                                                                                                                                                                                ?��W�  >�[UO >����0y���u�q�wK��6ՐR�V���\-|��Rv濚�Sʅ5V������P@����ŉz�"}簿6�%�0�z��@�'���"?ӈ���kƿu��TY@�6w�ۧ������*�����Z�^AK 0�ݴ?ې���f3@@������T�EG"A*����Ũ@W����Cd?�6���<�?Fc��o�*��k���?����ܭ��-��:ٿT���ٱ\��w�7���ъW���
kK�s��@���pb���5q|R��Q�#*=��@P�6L�?�u#]���6�PE�@�y��\��DB&�`[$��]��ÿ�gKב}����k\��n@�i?���AV�m�4�@s�5Gj�@D�!���=|ҙ_5�              @���H�5>������@���	| f@��8�%wA��xt   @�8`uR�N@���|�@V|�����@ ���
6�>s�6�w�?\݋�@?��ۗ'��D�     ?�<�^  B��dJ@���� ~{�$�U��o��j�������KB��g�û��!}?�����=�        =a%��nϚ?s��4�?<u"ʡ⥽�c��K��j\�H�ľ�� V`?QC{ƚ�-=�/�}>=�����?��a͖��@G���s�@�C(R��@ ���
>s��焼?��ۗ'�?\݋�@?�      @/��[W>�                                A�e��@  BL+��  BL��                           >܋���@��=Ğ>��z�@���8�=I>�?��m�@��Β��(                                                =�C U<@Ғ�x�?�7)H�+������:#�>TXqP<I'?Q����=�6���?�Ѣ���?;v�}��9�ث�-�=�)P�Ñ`?��t�G���h���4?���G����5׊#��>2�t�u_>k�롙����<�!1                                                                                                                                                <0�[B��>!9�S#`=����i��h�$7�Z<qB��u�=m��a!	<'�N���>9�M�1�P=��uX�滰�𬶃 <j16��=�噻S]�<-�k���@�i� !>��`ml���&�����!q܌�>t�
5!                                                                                                                                                �)�|�Z*>Â��!۽��>��ƿ��ơ+dȾ� �-^o�>glu�`DQ�(�I���>�dV!U�>6�,��>x!1tݏ��j�}5>�e���1|h`]f>/�6;��}��sf�R��8�ˉ�y����'>a�ىo!�1|`�?�f>/�PYK=�����0>
�VV��1|q�<�>-@bh}|`@&\%�G� >4+<�  ����˃�y���i�[�v�\"o��֑���@�8D�  >@8��` ?S��'?�w�V����r��]��(�3�                                                                                                                                                                                                                                                                                                �&1m�Ӏ >D�\%�� ���!K������+���&�E z��?g#WH�/G^� >J�0�i� ?S��,x?�w͸jZK��˾��p�]�גJ��@G\I����O��hm�T>�qm��J@��J.2>ď4�W_�>ՙb��F@K�흗
̾X���T�cy��e��w�Y�DA/�и�}�?v��O�Jq��ׄ�h��>4u�4E=�����QUI��@m��&�F�3�<�K�]=r𾷗��.><�����G�)ŷ���?�w�dB6S��$J��.'�_\iXf�z�bHޛBq�=o񓏝��=���׆�q?���[�a��)����}��?Y����",|-��>8�Ig�S|?S��C4?�w�P�}z@+[cK�v>P�jԪ��BX�S�Ͱ)=�fG��              @�i���ʾ�S�?@���	| f@��8�%wA��xt   @�8`uR�NA	X���z@V|�����@!3;����H��/��?�]2I.@8�	^~��BX�}�'���ȫJhFE ��O��[D�7��(Dzv�$��DO�wn�Di�IP7�C0N�b �?���3��        �����H>a�p7��f?L�`)�W��`��m�E=�%��W�UF�lئ>�y��:v=�� �lf��6om��>�����X����ɢ�iU�=�l@!3;����H����X~@8�	^~��?�]2I.?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?����O�
�=g��R�@:���$0fAnt��%��@:��TCAg�:$z�3                                                >4ED� *3��
ل"���v>"g�*=�)�ot�������]?��_�!V	>��;�L�%?�f�o�鸿R�fY�оA�� 6�����8A&�?�Yt)C!=۳�q�8�?�m��<�d�(���곟���V �?'�������K2;?@}                                                                                                                                                <Q2��seL���\�兜�����e,<o��і5#0=���lT�<�&���>/��V��Ȉ�z0߄����m�*����LQ>�~Z��R\|���X�)�O9�>�~
==Vv$��D#��I�3�>~����                                                                                                                                                ?�c>O���G�>"� fu?�;���3���u�s���Ǐ����-��P2mnݰ>kv���8�h���T�k�e mϿϚ�s�� >�������%8�k
p�>���i��d���I��.�?�n�U-���U�A;�!��޵S�3�蹌q>�(�ΕDI��-��?��_[Uy�3��&#?/19 ��`@!?	>W� >��0+�� >�f�"�v��˾���uGIٻp�S��yW��G.=\	��§,okӿ���9S�@��j�,��#��g�6�d�Z�                                                                                                                                                                                                                                                                                                ?��F��  >�+�?o@>�3�;����%W�����mD��U��ѩ&V�G�6�$
�§�������?_+@���'���#��.� �6���@��)��?���v:�b���t�@��Kā�����+�����X���6Aؘ�_~�?� }+�_@!�1�J�E���3a��A(<�LJ@Ub�~�r?�}A�@"?Ak���D��K,~�rW?{XX���-��jz�_��9~����
u*�}���tL��ެ`��@֬�f��j�ߤ�s�
�B� P�@I�`F�D>�v��ց���(`�k�@��;<)���},���M����
L�&��>���qa}]�?�S*�R[����y(^�A0��L>@*��*�b�@R� X/=����?�d              @�i¡�>���q@���	| f@��8�%wA��xt   @�8`uR�N@���80$-@V|�����@!2���>(�|��	?���,I?�Nr�2Z��R�    ?��5��  B���g�.@�K6IN��$���_����G�����uX����9{��?����G��        =aպ�xi?rF)H��h?=J�)2mP���=K������"(F�������?Q&p&�=�>l\���=���u��.?�L-Ʈ��@F�e  � @��͐�1q@!2���q>(���?�Nr�2Z�?���,I?�      @/��[W>�                                A�e��@  BL+��  BL��                           >��L�Ӣ�@�]ǵ�>��V���@���m�ؠ>����D�Z@��ܬ�;�                                                =�����0@���% �?ѻ���r��7�r��u>T]��x(�?Q���6�=�ʄ�(e�?Ë��Kj?<�{Ɉk�;s�R�ҕ=�/�h�Z?�#�ʖ	��9;��?Ȗ�3%�5�6/�>3�~��V�>k�����$� 	� \�                                                                                                                                                <��`'�
> �g�Z+~=��@��^���ʡ�Hb<qG6*��+=n]D�z��<(i{u[Z)>9d3p���=�?�#R[���,��<j9L�H�2=�>0�ɕo<.����+�@LT�J!v>��D-缪1�1�7��Q�*�>uCXl�                                                                                                                                                �����I�>�c<J��#����������)<�M�>gcY,�t���gR�X>�h�>5��LAY>w؝���+�5��#>�il\�K�1�	��l>0O �0�Ƈv���6����I�G<�y��Ȃ0&>av��b���1x��>0A���b=�?cK��>�iv� ��19�J&>-�a����@&\&M�  >4z�\� ���U������|ف�x�t`����Ꜧ��@��!s  >@��c�� ?SO,SE?���&t�.��p�B��]$|S�g                                                                                                                                                                                                                                                                                                 �$��B  >E@ʺ` ����1����bTB��]���:�֙pʛ���.Gg�  >K����  ?ST�+�?��݆�4���墿]$w���@F���ڪ�P���>������@���E�(>Ę|;�>���fS��@Ke�ƺ)|�X�>�P�c%�	������nȜA/��Dl?vPIUo�h���W��>4�_g�=�s����R��o=��]����0<�2�&%;ܾ�#�?Dp>=X�$�P �*�pӥ��?���Gz�{��:�[3�^�@a����bVĄq�*=p1�F��<=��"(չ�?��X�S����`~��h�֙be�@��"��8� �>9�jH1?SCa��P?���L�{�@��+��>Q���ݥB<�/����<�a�d�F              @���%yd����0,T@���	| f@��8�%wA��xt   @�8`uR�NA�<u�@V|�����@!n�"��B�y)���}?�n�U�n@?ѐ�Z�4B:�����B"�i%���EJdf<x�ϙa ���VG���D$*e;PNDs�h�Y:��_=0P�?���3��x        =�v,'>OBbF��?L�h$ח�=8����_�ě;����G�	Nv>ͤ�����Þ���=��'h�U�>����/���O,�2Ud�?��H���@!n�"��M�y)�f2'@?ѐ�Z�4?�n�U�n?�      @/��[W>�                                A�e��@  BL+��  BL��                           �э�?Is�=P�I��"�Jt�Ap�I+��n�#q��
ڰAju����                                                �q��J����Xt��Ƨ?Km�3dUX�)��d�S�p� ���?���Eˣ�h��ȹ�(?�W���Ƌ�Lǰ�*=�=ůΜ#>ǠA�$G�?���vޛ�>ij$�DH?�������"	�6���>ں��� �
��xu�X��E�6�f                                                                                                                                                ��{���=<��t/o�3=gEf�x��E��j����W����t=µ��^��$����>+��t|O0�±�w;b<ff�ޠ=>�w��>s3/����.=����&n!EHM'>��8�;��Q��*��d=��kd� �>z��ߕ�                                                                                                                                                ?��q������b��^�<|�ֈ��^Э�R����+F����8ݠ~1?�`��"p��b���S>5�0�! c�s��}?��T�"�,>�%�X�y��"O�:�!V�ֽI��&c>]�+��?��ą�����3�?4/��V�n�4\��>nb�ĥ7���}>���a%?�����>��4��T��?Y�B`��8@�F��  >�*��� >�Q�<"d���R[�|��p���U_jS�m��>K��?��nR�B�?�0]�	֪@؄��zz�=��!@ /aQ+_                                                                                                                                                                                                                                                                                                ?ϥ�H@  �Ҋ>� >�]E4�������JC�(��Rj���P^��,�P��ρ�?��R�0?�0`�P��@؄�
���=]C�+�@ 0.C�'�@ţ�s�����coD�6?7!&�YZ�@�N��p�@���?]��V�1�UA q��_�?�IY]��I1*�,����S��lA$���`S�s�,�]�Ͽ���F7�?K*=b����i��O=M�i�H�H+�7{�i�?��jd�s�Ƿ`�y@�����G@8^o��P@�!f��b��$rP��@r�Fw@B��fƼM>���܉i���4����@���c�������"�0˪�:���m���?�E��^!���N��{+�Ά��$�A�����
����@�+rɨ=I�q3�              @���u�>�P���ʿ@���	| f@��8�%wA��xt   @�8`uR�N@�8ےZ�"@V|�����@!nd � >!]�M?�?�*�pM?���R�N@�    ?z����  B���B�S�@��-���Y�$�.��e���SJ�����4G�O����z�Y�?��찁�        =a�Vn�:?qy���\j?>�f�ｧ�k�nya�����u�6��Z��?P�@,���=�M�Uy��=�8���?���t���@E���YMq@�1{wXa@!nd ��>!`U���?���R�N?�*�pM?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�6[p@�+I�CCp>�^��g�@�.�>���ӄ�6@����!�                                                =�w���1�@�è��?�F���r�҇r뼣>TgԀs8?R'�M�VD=�b/�f�M?�H�@��}?<��=<	��=R/�K2=�:wg�?&�X8�޽��A���?�<H��(I�5��aL>4��\RR�>lɘ� R�� E�&_�                                                                                                                                                <6�}!�> ����=�P����#��p��PrZ<qOL9���=nΩLm4�<).�N�	$>9�4�<�=��#�p�������<jF����=���.4�</�~;��@T���>����ټ�H�!x�����Q>u�w�_5                                                                                                                                                ����^>{����н�~������tľ�9fB/n�>f�@C�9���T��â>z�H3��>4�z��>w�3/�x���i&��>�۲�:��0�A�ܡJ>0d��߽Ơ��??C��evC�3��y�P���>aD��
%	�0�:k��>0d�t�#W=�Z��B�>�]�D6+�0������>.rW��Ix@&\&�M  >4�5K	  ��횃���fߎ>�a�y�Y�P��F�>�,@c���  >AEU}B� ?S(}��H?�nF�s��I�>���\É�"X�                                                                                                                                                                                                                                                                                                �#�R�n  >Ehb��  ���p&��h^A����S�ڥ�����l3In�-_A�}  >LF� �  ?S(��\?�nFm&m�J�H)�\ÅX{�@Fʁ<L�PZ��3[�>�$Z6��:@�k.%���>Ī݋�2�>�T��T�@J�Ȁ�f�Yxʒ��c'��t��nq����A.JSB?v	���&�����>5�*kNz=�L�ͳ�T�R�LI(b���Sv�<����<���������;>>��å־+o�Ժ��?�nHD.����]?�!���^��P#�bm-��+�=q����M�=�K}F�0?�e��f���_�̊����.b�G�#T���>;{8��%?S(�
1F?�n+5ǚr@S���>R[W���2B�!�/���=�u�T�+              @��c�=տ�?��~@���	| f@��8�%wA��xt   @�8`uR�NAz��m��@V|�����@!��AM,_�A��t��?���/�@G��$�;�Be���P��ejP�'E94uWk���@O���78���sEW���8D�d!��*jC��p(��?���3�K�        =X!2�)iN>(�c����?L�m͔7�=�|��x��J�7)%�+�?���>�Ϧ��NV�Q
��=��4�>�'�81�x�6�XAl7�?�J�zE�@!��AM,t�A��t�<�@G��$�;�?���/�?�      @/��[W>�                                A�e��@  BL+��  BL��                           ��>܁����8p���~�@�˔.Y�Aq�=��s\��dH�բ�Aj����/                                                �;���9��18a��?oXAއ/^��r3t��`?A��a`$?��tA�]2��tE�ŪF?�l4�ҿB��6�>r��?�@�ȇ�
?�i��#�>Ǖ`~�D?�l2��Q��� AL݃?,�qk~zڿac��O���>_ftY                                                                                                                                                �W�������y��F�=���q�<�#Lsͬ=]�qm��=ѷ����=+�ao`d>#��"A�ؽ�N74�<�����>��Y�>-2�8�ƽ?Ce�Ǌ^�϶���>���^-�u��'-�;8=�L� ��>r�EHi(�                                                                                                                                                ?�ꦶ���M��Y�.��� ��s��Zq،32��m�J�2U?S}I�Y��@v�vƦJ���c��z=�_��9z��_4��V�@j�)���� *�����~�#�.�aҴq%q>���ɆLB?�qY�x���"�P�(}?��#�$7|�5սA�`y�`����?F�%��Į?p�3�`��;Q����@pč+F@=��  >��$   ?��������ysk�k}h���7�M�UN]u���%!A/tH�/�.\���@:tm�!v~@ׯ�>�;��O�W��~@p���                                                                                                                                                                                                                                                                                                ?��;X   �hug
s  ?���	*��yr��¸�#Q¼D�?����E�r�%�xG|�/���@:t�?��@ׯ��nel�P�ys�j@pV��U��@���'�Q����˝�?��@�@y�l«��@��Qi�
��4����A����-/���\s�������i%���5l.R�A!��;�ԫ����~~�#D�@��F~�s�bZ�<��B�o�G�f��)�i�Iѳ@*6�(�%����p�
�@t2`����@�����
�@��Y8����tU��$@��r8�@6�4�%�?q��Q]-���fv�!a@�M��@!Ja��A��u����A	�����W@+����̃�Hӏ�����8�k��'AS+���s&~ރ��A�^;����=��RV�              @���EEž�F)�4�B@���	| f@��8�%wA��xt   @�8`uR�N@�k��cS@V|�����@!��5���Q�Z���M?��{'�V�@'y�R����JT A��Y[�>Du�4Dc�B�ɗ���r}�|9vwCT�t�ˡu�$2�J�z»�*gw
y?���3�<#        =����q2>���k(�?L�K�W=�Gwqr��O��w;��p�����O>��[�ʫ��X'Z��=�_^��?��g���?�q��k?�{�١�@!��5����Q�T�21@'y�R�?��{'�V�?�      @/��[W>�                                A�e��@  BL+��  BL��                           ��^ �x���X�#��9�?�e��0�Ak��v�BQ���x�.'A[��$=                                                ��=1֯�i�o6P���ǴQ0]�>$��T!1���ȁ]�?�△f�>/\��s?��@�t�?]T�D�g=�y���>h�L�]��?+Ȁ�$;\=�|�����?�T"�1�2���o3>�7{q�����ԟ7�f��Sy|p�d                                                                                                                                                ����1<\ƾ+��	�`a��*��88<A�U׈�J��Y6p�t?=⭋r͞<�4'@k>?�#8S=��%&�<O�a�'�<�'��@]�=�^Ζ��`;��z�0 #.��>���+��?�)yxu#H=.C����>��m���9                                                                                                                                                @".,8j����OtZ/>2/3��?�8y�G��؂N��R�����>d�:@���`�6���`��2���.�6��?mڴ��}@U��nޞ>߆=�&�4B��gh�>�~��gr�>E����2����Y,]��DN��a >�ٓ� �1;ËYQk>�.!�s��>g]Y���[?7�����1;%�,Å��yc4�l{@%7�� >��8�� >�.pjA����s�jӿX��پ���F!R3Q/��i�@�4?p�.��M?�;�@�ifxa��eK���3?�2�E�й                                                                                                                                                                                                                                                                                                ?���*�  >�2��� >�=�ג��p�u�����D�F82��t��j��7�?p�2�L#�?�r��@�ig~�"��e�_���?�2��%@��d�Tx? 7�aLx�+<���@�!E���A��n��?2m3o��lA���v�쿍�Z�>��D��~��ٟ�-�EjA+��E��;)S)?��#ZS>����5�:>J�`�~�������п�c&Zf�l�Ů$q>c`�x�,�`��?w~A���?��̭*P@�ր��K4��gB�i�@ �bnxP<�:��K.��Hx��ʾ�Gy	�@}6�z?��{�SɿC�����vLy)�?}�F҃�?�<��W@�%9���@�~@��J��M�V|��AU������<�As ��              @�
i�7'>tT)r�5@���	| f@��8�%wA��xt   @�8`uR�N@�⊑p��@V|�����@!�VA"�=������?udRX@��S8AE��|�  �R櫇6	�D9�k��B����Un�E'��c�?B��7��"YC��(w���BY��s��?���3�˹        =+�	�>��� �3J?L������E��=-Ǽ�0��V�@���/��U>��%���=����<��=�<��ǉ-?$�Iאȿ�\P��6?�
���	@!�VA"�=����6ͺ@��S8?udRX?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?��Q��Ż�=^?b�윈AWjI_^�?�M_�x��AM�y��                                                >�~ƈ�Z��t�D]��	U��վ]JO_D��#����?����u�=�}��n/?��0O _?R���=t�^�hd�>U\̲֙�?!�.��ܛ�wg}=3s?�u���)�4Y�]ð�>�p�K6�>�CJ# ����ࢄ�                                                                                                                                                <��:^Z� ���t�6�h�k�x٥��M���X��=�[䠁X�<;q��Ae>9މ��Vc=ȎNV��9����ys�<����X��=�x	�zY;��Sĭ&�0�#lL>��a�����f�e�*�B��]3�y>��|���<                                                                                                                                                @�a��c>��[��;pu��p��@��x픧��	Lw�+4��F�4N�C�"���>u=���\V���o�Dr?�'��1!�=�Q��:����~h6��0�� ]4>%W)�W�L���gސ����(>�=(�&R>�5�3���0[�6#%�>#�(�bo>Q-�Eeh?>�iM6�8�0[�{F���Q&"o�Uh@& >jp� >�8A6+��Y��������"K�*�;(��O�7��dL�����@
n�?B�k`?��h$�@��[Λ����lS�+��0�!��                                                                                                                                                                                                                                                                                                ?��b��  >�w�xXՠ�vܴ]��������'�-��%b�˿7��,����ѤSV�`?B�R;��]?�� ���@��v�h	����῏1���M@������>��X��9޾ؼ9��	�@����n�3�*P�S%5���YINtx @��cP�(t�\t�igb̿�%E�f�i���:��\�A,��m�'	���Z8~�w?�F�$�gn>�1��g%f�n�Hs���?b-��+n��1��<پL�RP����=	g&!6�?CC�[��?T���#@��*��F���U�Y5?�Ь.)q�@:��P��g>��ȡGT�>pC�p^@bP���{���u^�w1�7�*9d���*����?RT�ϡ�	?��t���@������@���ĝ\?EZ^�V�t@!5T��[=W/��è              @���o��>���E��@���	| f@��8�%wA��xt   @�8`uR�N@��E���@V|�����@!��U9?>#K.�\?⓼^�?���zN�@!5     �� !��  B��~�w�F@�D2�����%��������*�������5{��s��c?���O�n�        =ae��?p�2�H�?>�+�qch��l/i�㞼�:�:� ���2���?P���4/=�\��h�=���x�u�?�2���q@D������@�d��+�@!��U?�>##|lf?���zN�?⓼^�?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�S��4@�?s�&#�>�!�,�=@��v�>�K�F�6�@���1i                                                =��{�9@G0d{?�ٽ�6C���[A�y
>Tt�x
տ?RiM��]k=��[��?�	|f��?==Ɩ�G�?:b�k�=�H�~�*#?hQHg;㽸�3oM"�?��.K+|+�5�)�#,>5{XQt��>m��&�p� �}I_ћ                                                                                                                                                <��~�> Z���=엥�O�����v�T�Z<q[�ZnG=o=�uc><)�[X��>8�I;�=��~V�O���H���d<jZ!<� �=���Q��<0E�J�&��?���u��>���3O��z)*_�f�����I>u�(�e�                                                                                                                                                �X��i]>ݹ��hf��=v�ϐ��Y�4����P����>f���F���Xf��W�>�o��9>4�ߡ,�>wq>���y�9��=�>7m:�(�0"%Rh>0�[��ۀ�ƾ���N`��=���؅�y�鉶�Z>a	r̬��0"��j>0�L�7��=���G
m>�.���S�0!�����>/E�	�"@&\'l-� >5"��� ���;o����*g�B���{�D|�צ���P@Û��  >A�c88  ?S6��J7�?��S�N2b���9���\mc��@                                                                                                                                                                                                                                                                                                �"���+� >EŲ"X  �����1���+ףD)꾧�U��:��W��k}�,��I�� >M���� ?S6�M���?��T),���OӖ��\m^9���@E���u��P���U��>���=23@�.��o�x>��8��iR>ֶ�!EJ@J��\����ZD��k�c6�b�6����i�!A-�T�n�?u�E'�����>�{�
�>5j��=�*��Q��S�E�������UT�g~<�@n6҂��r�[zy>>��XNe�,^�9���?��V�Y�ߍ��vz�^Ro��꽿b���u �=s�/��=�̃`��?�4��w)پ��}������Wo޶��#��2=�>=�#0p?S6��nE�?��6���@�����)>S87��L�Bt��~=$����              @�hw9d�i�,*N ��n@���	| f@��8�%wA��xt   @�8`uR�N@���Xy��@V|�����@!�@%�����-��=?��tmp:�@.�E���{A�oD� �r���>D� �!Ǘ�ët���LDx#n��r,D
�
���T.��<�{�J�,x�?���3��        =�[gl�>��I5t?L�>T�Y�<��n���*�����g?q /2�>䈨����=ǻ9�N��=�>�:G��?
���?z�mxwn�����@!�@%��������@.�E���{?��tmp:�?�      @/��[W>�                                A�e��@  BL+��  BL��                           @V5�R6�t�pS
�O���V��NAy��ׯ�?ٸ~i봿Aa��l��                                                ?�E��K� ����I?��?��a>�#�Mi�W�B�4�\?�����ƺ��+7�%GE?�J�c~/3?m� ��	C>_+��د>��@��c�?pEVk�'>*")=��-?���=<�&�1e�J9>� 2�*�>�R��,���
��O�t                                                                                                                                                =#O�\gξ<?@t�o=�{��ޠ�<�-V�#;�_����wp>Ϡ��H��"�phW�>Fw�-�=�z�LA��<�?��B] =$�{g�z=�#ObUס��R`́�|�/A����>��X��=t�-*G�٨�HI�zkJF>���PWV                                                                                                                                                @2-���*?Jj���>�������U�U}~m�V#�r�Tsr�@6^�i"?"� .��">�/@������b�U�@8l��Ap�?�:ԓ�e(�<���¿���[��>�0A�׷���m�3��+���2?pj���`�2hn�!����#�	�(>�����'?��|�,��2s����?$r]����@$�(� >��~X�  ?�Y�.|���vZN��dP��2[�K�^�r���\����?S�X���0?��r=x�@ÊT�zJ9�R��+�Q?ٲ(-��                                                                                                                                                                                                                                                                                                ?Լ���  >�w���� ?J'���*�����n��Z��6��`FM;*\��զ�?VN\��?��F�+�!@ÊLm�fJ�R�	��?�6q~��@�A�`������Kܿ?�M���}@��Z\�����I�Y����;VA����?�@na�ɜ?�*����߭����A)�����@8	���F?��k��#?lhK;�N>��/`�Z���։=
!��oȦ��$~DuҎ��t\n=�N?UyX-��0��)}�$��@��x/c���Z"����"8�����W�V���NcP�!�؏�c��@�}c6���@�^C��?]tU%���J�[���?]?u2`z:?�"��c@�{qD��P@�H�4.�����d|z�Ak�%H�<���ř��              @�h&<4�]�����NV�@���	| f@��8�%wA��xt   @�8`uR�N@�F��sqs@V|�����@!�L1����#��D�?m�Y�jș@�Z��[��k���  A)5�Q��D0�T�p�B���J[�(g����B�Z��D~C���i[BZ���6��?���3���        =&v�j>���2��?L�^r!*�S����@՚i�ξ�o���?X�I��8=��d/��=�N��[2#?-����]ÿ��DAQ ?�<c$Y�@!�L1���� �{7R@�Z��[�?m�Y�jș?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?�N�� ��0h��E���IL�=�Q'AN��8�?��jr�fAD�����                                                >�a�
;a��[=��f���h�$W�j.��*�!��~3��?�F��=�ͽ���^���?�*���n�?Q}"�bT�=N}�D�&�>L���0�?!�}�Ӱ=�
z��+9?��M�B��4��t ��>��=�~
�>�  �]S��˳�O-                                                                                                                                                <��A�Ţ���d��]�EB$�����6����̼�,e�˘=Ԙ����ﮌf�x>8�X��`=Ƹ`#O|�;��D\���<�4S�V�=�=�G�%�.�D�.O�1?���p�>�mڌ]���X��>��+rj�>��̦��=                                                                                                                                                @gA��>������}(3V?=@<@�s)���.pt�>��%9� ��	ZOT51�>p�8M�R���N�?b~�?��������v��;>�Fol�B�0�!09w�7�o��=�/�97�~��?N�p�j�(���D}+>�m��Q�/�"��X�7���?>Ea�<r_[>�0��hu�/��2 ��Ru�A*�@&0��  >��c�� >���W)�*����Z��*,T�]�ǿ00t9@�o�¯�6R} ?'֧�o�a?��gW>i@��b��ߓ�t!������Kj�                                                                                                                                                                                                                                                                                                ?�qB��  >���Y� >�@�}����=Ґf���7J��08+�|
�¸~��E@?'ؔ�ӌH?��5���@��	�ֆ��tn㢅�����}�@�N�,ɩ?!]���ƕ�Yԓ�l@��^k�Qߔ2ˁ�K
�g@�?���I��@�!#�A����}fwX��bh�]�A,}�k|��?��Cz��$?�����>�Yz�Q���3�g�?�������p P����#���\M��r)?(Uc6��Ͽ>�ОM@�ݸ)t����&>a_?]Q�؊�@N=��0�U>��S�B������G.�@V;�[���8�<�g;�1~$h6s��h��A|�?7u.1�Զ?���N,I�@��sI�0@»��M�?U+�%���@I`��=��d��s<              @�n|�H�z>�|Ӵϊ@���	| f@��8�%wA��xt   @�8`uR�N@�i��.\@V|�����@!��X��1>_t#�~?�	֡�?�r����I`�    ��ʽ/p  B��]�v@��Dj�|�%g%�,����Wr�Ѯ��<� ��R��3�?���k�        =`��?o��&?��??憫�h�����ּ�F�f���-ʶ̟C?P;p+�^W=�n�+�X=���+^?�W��۾@Cu � �@��i�t��@!��X���>_o�p�"?�r���?�	֡�?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�8��@�_,��Y>�s)�1��@�6�.L�? ����@�#���Fh                                                =��>��
@��f&�V?�a�!�~ؽ�@b�>z�>T��d�??R��Um@f=��	���W?�§�#@�?=�h�����@��i3=�_��Vc?���E	f��o��i�?ǅ� ��5��c>6��#GpH>n��;�(� ����                                                                                                                                                <dA����> ����f=��ؓ�~��UKg���<qm��`�C=o���!H<*�:H9ʫ>8_D���=�d<�ܷ廵��47C<jw��@�G=�Kʃ��<0ۧ�a�+�?.�R��F>���߉����i��Y��c�C�D>v9��mN�                                                                                                                                                ��S:\,l>V�����i�B�L��₇��h��v[�r�>fcevnq�����p�>T��Uo>3��
V>wL���<�v�����>­�6��/U�m���>1Wc�t����M��9����I: ��z�"Sn>`�%��[?�/U��2^?>1GsVbw=�;iq���>vx;��Z�/UjK�CH>/�U�f�B@&\(A� >5��[x@ ��Z"1������9���|�I�҄����Z4�@��8�  >B�{R  ?SMP��k?ݫH����Y��	�\��fؾ                                                                                                                                                                                                                                                                                                �!Vf�� >F8>@�@ ��^ƥNy0���/Z3u���U�!�3_���S�=�:�+�l�  >N?�H  ?SMVC�?ݫ�����<z��ǿ\���JO@DꑰK��P�����>�i��N��@��s�0�>���tKDw>�.��!0�@J^����[E�I:�cM �׷����`uA,�Az%x�?u��p��A�|��1>5�޲���=�+/���Tڢfv��U����8<�u���#���AIn>?�C�q���-��0�9?ݫ�����׶vv˿^����b�9no-=v��]&�=�����?�6"ĸ�V��Y#�Bھ��B�ח��$�-��Ɖ>?1WM��?SMA �6�?ݫ�����@���j�>TP��i�R@D���Aq:={D_���]              @��dD��">�
�0!�@���	| f@��8�%wA��xt   @�8`uR�N@�t~��@V|�����@"!��ܴ�>uȣF��?z� �&m?�'�;�K@D��    ���2�
  B����~�@���6�a�%�q"9���b�\����v�T����_�c�?���et�.        =`�3]��?nL��T�?@Y�/C�[����B����+20����<�?O�T���F=�}W�/Q=�%!pr�f?�Ņ<th@B}f?5�@� 9��P	@"!���Ӯ>u��6W?�'�;�K?z� �&m?�      @/��[W>�                                A�e��@  BL+��  BL��                           >���0��@݀�$}��>����p:�@�Q�l �?Q����d@�<�ڠ>                                                =��"��@��~�S?����ZJ�Ӛ6J�>T��	D?R��[�
�=�]�z�$?ߏޯ�?>V9���b�A�4�na=�weO|�a?��:�	��5K�ߔ�?�8��>¢�5٨��>7��_���>o�*.���� ��{�                                                                                                                                                <�X�X	>ղF�^=�*�AtH���s
�<q�d�?�=p�J�pf<+��&�$Y>8�37=�����軷M��#x<j��h��=����ÒM<1_��ۗ�>�gm�V�>��/I$Ｏ1{/�����$��>v��Md�                                                                                                                                                �;�C>�_}�%�7��^����H=%���OSv�>f8�n}L�:|�նw>����x>3���k�a>w;Z5%��j��>6��{�\�.�L�� �>1a�N��������:�� ��zQ�Qm�J>`��{<��.�=��.;>1a��l�=���VA>keA[
��.��ڋO>0=��T@&\(�-  >5����  ���,�b�����:-�~�a�7�վ؃H�	�$@HO(j  >C:
�~  ?Sd�
"�?�O[P-�U��jͭ1�[�?(7�                                                                                                                                                                                                                                                                                                � Z�M�� >F��I�� ����[O������t�˾�������5;Q���+T��  >N⻽�� ?Sd�,�Sr?�O[�0������I��[�:\��@Dk�>��@�QG��(�>�?��#@��h�"�>� ��)�>ח�8�@IǇ0Ⱦ\-�x�\޿cdo��m���O�����A+���[�&?u]��%[��no�x>6.�eȧ�=�	���?�U�Ωh�Ͼ�������<�@�m�)6��j��$>@WU���.��ƅZ?�O]�%Y��iW�ƚ�]͑SoXF�b�N�=v-��}^=�F��B?����W^�������5(���6�%pk�`>@�`��R?Sd��~��?�O8�8�*@oC��Fk>UPF峈�B7�ZN�.=�"$�%�              @����n��
��P |@���	| f@��8�%wA��xt   @�8`uR�N@�P���@V|�����@"]���a��O�5� ?�� G�i@.W6e�"�j�{��B6���>eCD�Dz�$�#Dڜ�DBD��hY�"ND�K�*=�)DT 8�>�C����"�?���3�P        =�#�'�,�>�9�a�L?L�<$?̽�l�����4��` �g� SH�k>�s���>j���Ţ=�S�9@ ?
�@K��T�Yx��Z��nr�@"]���aɿO�5��@.W6e�"?�� G�i?�      @/��[W>�                                A�e��@  BL+��  BL��                           �����AmABI���w�@��{�`A\٬n��*@M%�/�Y�Aa<�	Ȍ                                                ��+���iK?�/��*������i	w�(�Q�%(�V/�����?��ixw�K?2�.��?�p��ۿg4�!	h��&o�d�I���w}��!?�7�mѣ>�KIؐ�?�J� ���1)��|�q��7�iJ�?6��k�G��	�y 7R�                                                                                                                                                ��Z�q�n>�5����צ��]���D����r���8�=��Q�B��=���<]�>*#�:��%�Y_�ѽ^4���h��x��>���ߐ�[:��_�0��+�>��[��=c]�Ѿ����K-uy�>�6U?%(                                                                                                                                                ���Ao���J0����;����?ͩ�ˎ8�ӂ��Dbp�g�h����� ϣ�M�6��K𔰏�?�(?��ҿtsl�D�� ��d�'��������?� b����p?�(�O�3��T>�p>�Q?��kM����ǰs�l��*~Ɨ�{�/1�za_�NLY+�4���<�k{?��Y&A��.����ڠ?�PFH�Q@$1�� >��r�   ?��6x����i��9*Ϳc��I"F��J\a�c�D���+���5�	[���3#V�@�z�#�0Y�(F}�MS�T��;�H�                                                                                                                                                                                                                                                                                                ?ӣ՗p  ?h�ޢ  ?��%.%����g��K�u�
n�L��9�(&L���{1 M �5z�X4���G\�!@�z�F8'��(�u ���T/�ɝ!(@�|��8F@�I���?���Q���@�v_*ğA��i:9�%��N��hA	gi�]�\@�y�>�����@[��o��ᎸQ|!�A(ea H=@��)��@\���@/J�?/���C�i<�\?�?��N��@!�	�z���8Ό�����<s�?�yW�-�d�
l�x�),@���WY%���As�]���Ÿ�$@[�A�I?��.�$�v���r�`@�Ck��S��<DR�O���0�.�?����K�7�@�A8:*�� 6>�ޱ�@������@��_��@A�.-@[m�tn/=�f�\.              @��g��[>��c>�@���	| f@��8�%wA��xt   @�8`uR�N@�� ��ɘ@V|�����@"`�G%Y}>��??>�ʇ �?�X���0�[m�    ?�5lJ�  B���\�@���+��&#S�B��^Y�� ����S���z��FG�� �?����w��        =`���ъ4?l��_/��?@�U��	콦Nl2�u�����vB����1�?O]�e��=���~�6�=�z��r��?��慃�@Ab��ӻ@�!�y`�@"`�G%	�>�;Zn?�X���0?>�ʇ �?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�T9<Ş@ݯ�$%��>�!��;�@�wK�]چ?N��M��@�a�                                                =�T��a�m@�.` W-?�3���`��	J���^>T���I�?S:��ۈ�=�%F	�{z?�JK��'?>�o���B�"O!$=���Z��i?9���$��"��}1?�������5ٵ��K>8�F0>pl��r�m�<[o��                                                                                                                                                <�c7�� >f&D�]-=�x�׬���������<q�B�1\=pPd��´<,���_>7����7�=����u⻸�=C�k�<j�P�.<=���O�<1�w�]z�>U�H�V>��@t����]�G �G���ͭBz>v��6Q�                                                                                                                                                ����&)>B��苋��ԯ�W4��$v#����sq�:>fz�y/���hR[>AFk~:�>35����>w5{�J"��sF�4�G>�IN���-�̨�/�>1�����D��7]T���@��ܾz�Y��ӻ>`�N�t��-Ƚ�yD>1���W�q=�~�z�>i������-�\8��>0�6a��@&\)H  >6Yc8� ���0N�*���s�n�w��]JV�*P��8UR�@h�  >D�jh  ?S�1��5�?� 7�lC�>��e1��[���T�                                                                                                                                                                                                                                                                                                ���A  >G��� ����	ԗ��u8�@օ��C�J7E�ش�­�Q�*l98�� >O�I��� ?S�6�~k�?� 8X��>��dSA�[��H��o@C��v�<��Q��BL�^>���L��@�w�_��>�ct�H<�>�S7Γ@Is�Q��]RPϙܿc����7��� l��n�A+?�^L�?u0 �#�T��u(����>6����d=��XI��V�t9�_߾�C��ľ<���D�Ҿ��k�u��>@�_�]0�0
��6��?� :m�x���H�T��7�]��*��c0�F^`�=v�.M���=��
c���?�:�4Ԇ��F�S���ش��&�u�&P�����>A�˶�R?S����?� ��.@O����(>V��]ԶfB._����=Ջ*:              @�f�����nMt�Զ@���	| f@��8�%wA��xt   @�8`uR�NAz`S}�W@V|�����@"��P��n��YF�7�?�l��d-�@3�Ӷ�t�Q��/�B,:�/��D�����Dr/P�uT`D���\9�~Dl�q.?�DU��.��CMk��d$?���3��l        =%�vR��>r�Cǟ/�?L�SL��H�g+������j���� �`[��~>�貳)�=�L��=c}w�:N ?N��x�=�_��?��!���
x�#�@"��P��]��YF���@3�Ӷ�t?�l��d-�?�      @/��[W>�                                A�e��@  BL+��  BL��                           �Dpd�NB��Q�
Bd@F�2y��Ag�1S"��@�G��7AdϪ�b��                                                ��E:Y���~�r�����}�ͣ���q�j߾��W�1?�g��5>�|��m`?���k�UyM��S-�PIf��퉿g�"[�?��7.`o�>j)���?���K�[�.*�Z���>���{;/?u�'[��͊ �M�                                                                                                                                                �M�[����+�Eg(���}�2D-��%`7h�w����Pɜ�=��8
�AL=��Jm�>0���Ȝ��崸45��(�17L���s�?*l>����0����Sо.��8|�	>����7����@�{b��\�>��g:	�                                                                                                                                                ?�6�()n �S�����FR�{�?�٩r.�<����B�2��8�������r�\0��J�ϾuI�얘�n�h�(��Ͳ�vxd���M�YS�$�]�G�??Pz�\���[�?�Gb�}�����*�������O��/�8�Ӟ]��9�[8�.�t�;�s?��
��qw�/?Vtb*?��V���@"��ܑ  >���H  ?L9z^��U���gH#�f�mמc0¿Od��j�K����������V?�d2��w�@Ȑ��`2�ݠ��p�`ͩ0e�                                                                                                                                                                                                                                                                                                ?ѪQP  >�:W�� ?L!0��-���m�i�ÿ���cS����t�B���f���
�F8�?�&<�܈0@Ȑ�0�"���P
M��;���@̽}�r�@W�q��!�� !abB�@�aI��������6pf�c���A�R��w@+�ѐA����#('���ݸ�ˀA&o�Yԭ@q��.��@l�D�9�?��e���Կg�<�p�]?�~�t\��ڇ�*�@�ʶI}�������d�ֿ� �8�bk���d`�@ɟ�6�~t��lN��As����@M�K�9�?BU�!�j7�BȘ���5@�LI�-��"#<�#æ����k������N�ʛ��C�c?wSWcV_�@��r��.A�?����?��"I�=�@O�(=�d=����Q�              @�l�&��>�s����@���	| f@��8�%wA��xt   @�8`uR�N@�w' A�@V|�����@"��&�˧>.P.56?��s��?��2��J��O�(    ?�p7��  B�R`�(�w@�������&�.��R���{�K�D�����w>e���t4��`??���#/
9        =`�)�+ʞ?k6���o?AF�Y{����(��%4��^ʈ�P̾��l;�l?N� l'�=�����Y�=�˧=��?�~��!G@@R�#��@�;Z82�@"��&��(>.SިXy?��2��J�?��s��?�      @/��[W>�                                A�e��@  BL+��  BL��                           >��Q���@��3ծ�>���M��@�����gH?Za�ł�@����S�z                                                =�)����@C9�<�/?�p[���_��}6V��>T��9��?S�B�(�f=�����o?�R-DƏ??^B����D?+�b=���A��?"��Y^���R-\?ƐK��e�5ٝ���>9�,�ٛj>q�E��c�zo�p�                                                                                                                                                <Yif�;e>�;�!�=��帻�b�W�;<q��m�=p�|��f$<-��Q�O�>7t����Y=�`,DF'��M�[7-�<j��=��=�T �\/e<2�����=�K�Q��>�� �{���)J�eV���->w+��I�                                                                                                                                                �-��s>��y�p��������|�E�*��S�ц>e��6���-A|S�>�X��>2ە]�>�>w?�Jl������>W~)���-��C
>20O�E�j����H�;����ށ�{m��f>`���Z�-���x�>20<�9#=�-K�=Z>s�i�!�-E��M>1�~tz@&\)�p  >6ϵe(� ��s �d�*��:� �s���~Eh�V��ن��8�(@yw)J  >D�C`  ?S�%�:��?�W�����$߱P�[_|�w                                                                                                                                                                                                                                                                                                ����  >G�a�t� ��w�RhuS��;��ZP���2"�b��9|�v\�)���� >P�xf�� ?S�*�2J�?�Wưd���m����[_ws	�@C]��O[Y�R	�Va&>�������@�>/�	��>Ų�>>؝�gA�@I,�$�ۺ�^�V��c��j1��� s�:�|A*�r��?u֭�D;��|nc�E�>7r���=�$?�;�XB�6�տ���2*XG�<͢�B@��L�t>��>AxG��(�0��[�0�?�Y��0���"d�]pt�8L%�c�9�z��=w��%Y=��\ �.?�iq�a������@�n��9f��)B�'?F37\V>C��Q��?S�ю�?�B�!�3@>n�)�>W���覨B@�n��h/=
EG��]�              @��h�z���WO@���	| f@��8�%wA��xt   @�8`uR�NAb+uF�t@V|�����@"�P60���u�m�Z�?�_=���@7�}�ڏB@ŘȤ�HA�f#��x&D�]bzRC�ɬ�U�D�T�|wշC�e��D]y��WC ��F�=�?���3�!�        ���髴�>eA��>%�?L�^�$�/�Y�aV:<��J���V��F��>�nx��fM=��+�}&$��J����>�d�����[(�o�Z����#�L@"�P60��u�m�巇@7�}�ڏ?�_=���?�      @/��[W>�                                A�e��@  BL+��  BL��                           ������B��1�u�E$@.@V0��Al��g&(@-��8@�Ag��t���                                                �x6�$-�������~濗 �{��*D� Aʹ���Bx�#?���Y�?>|B�'dB?����Խ�O������Ǖ���9�Ģ��?�s�E5�K>�Ѻ���?�����6�)�;H�оΞ_�+�Q?�GS)n���md                                                                                                                                                �����ݽ� ڟJ�Ž����<�3�FIL�'������4=��]*��<�[W���>0�_L��K��xe��X伐����:���wZ>	Es$3���ZA�7)�,��s9� >���B�=DKp'�C���9��>|�7�~[O                                                                                                                                                ?�Z]cx���z�j�=OJ4
��?����<�俳Y'|cg���f��X}� Z1��A����=�u�x+������f���� [�?�S���h5�}��$�A����>�'5�h ��3�v?���h�����oD��0m�����0A��?�>��m�|�̪:�n8�?����)7�0ECA��?D*,;��u@!��^P  >�lbZT� >�q~������!�-�tM٧���Q�ܡ�"5�������N�,����Ɉ��܃@�}�<�����J��>�(`��MM�                                                                                                                                                                                                                                                                                                ?ϗ~�@  >�P�N�� >�4���Q�����n���*a�E�U��l�
��Cd<߿��&5�����ɗg���@�}�z%���X�N��(`H\��@�X�'6��?�\��j�9�d�F@�@��t�D�(��#�SpsB�ޫ���89AOtP�=8?��C��@�k��p���w���A$8��=׽@U��}㡵?�L4l5�P?;�����ܾ�9Z38�?�s�&�(g���;���NDC��p����u�ѠZ��%Aɫ����7{�x@�<zEAj���ET��)7�Nd�x�c@F��M)�>��*���S���<1i��@�1}� �(E⭽��VW��52���re����zs��uk���8P�@z3[2�Af��l.@@Vb߼�@F'k$��=zf��mg              @��U!U�(>�y����@���	| f@��8�%wA��xt   @�8`uR�N@� �X��p@V|�����@"�� ��>�b���s?�WR�7?�͗�.�@F'    ?�9{�  B��u�r�#@�W�~O|Y�'<�1����L��M����A�߸���A�$�?���N� �        =`r���?i��zl?A�F��Q����)N�O��"�������%t?N)���D=����*�=�@�+l\?��~��8&@>�j�r@�O� ޤ@"�� ��>�n���?�͗�.�?�WR�7?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�8Zǲ��@�'�W2,v>�QgE�@��ٙ|�B?v����k@���.�)                                                =���k��@��?ͺ�:�	����z~�̮>UP.��?S���A=���D�C?���Nڵ??Ա&�u�E�#&r3�=��)rۣ?«�+^=��3I�J}?�C'A�B�5�bKf>; ���;�>q�W�r����o                                                                                                                                                <��<Z�>�����S=�8���������/2��<q�ɬ,N�=p��{m<.��c^3>7+�
N�=����u���߳�<k.��9�t=���Nz\<3H(ԾZ��=���8�>��ќ����	�p[i��\l�L��>w{����                                                                                                                                                ���,�>YB����6El��G���"�#�J��fʐ���>e�AφO���y�#7>W���r>2�c�i��>wZTe=��~~y�n�>딱��K�,Q�Nw�>2����\����ȅ+�� ?n�ʾ{�.GPw�>`���?"'�,Q����u>2��r�
=���w>�
P�,Q�e>a�>1~�B�@&\)��  >7J�UE� ��:�P��.����NV�����:�f��p�S�)@{��<  >E�fT�� ?S�w2k�_?�{�����ǘ=��[6ҾҶ�                                                                                                                                                                                                                                                                                                ����m  >Hx�]  ��?���aS���Ҥ����{�Ht:��ê��IE�)n?��  >Q2%�� ?S�|���?�{�B�j$������[6�0u��@B�i�]7��Rq#��ǭ>�J�^�, @��A�>��F!g@>�(�y�Z@H�'!���_�j�5YN�c�<�&x�� {��\A)��!+�?t�v(�3�������b>7�a��=�6��F�Y��������{�@�<ε�Ww}z����4��)>B�
Ə�1�0U]c�?�{ʙb�����?o	��]TA�\}�cݳ遢=y �gL%=��eLoD�?�����n�����7��Ó�r��(=g��>D�=j%?S�`8	U?�{�!6s�@;�j(W>Yu���'7BOF@̣=O�z��!              @�6��Me��p���*�@���	| f@��8�%wA��xt   @�8`uR�NA���$�@V|�����@#8��.�`��G�5?������@=���.JBOF7�J:A�ȍ�7E�+��C�n@w\*Ē���D�D�i�,�De���Fe~C'�=o-P�?���3��}        ���m4��>U�ٕ[�?L�f�d�z�T%�ca�=P��ݺc�K��@7�X>ͥ6��br=�ĭQ��v����~��>� ��

�R��lF)?~�Ϭ�9@#8��c�`��|��>@=���.J?������?�      @/��[W>�                                A�e��@  BL+��  BL��                           ��,����Y�5�NHR_�@77zp�;�Ap-r�q@7/d���Aj!bi���                                                �C)v���شLG1䘿}�[�޺���W������{$���?�+R�9k�>�;A�4��?���<�b��I�L��������G;Ⱦ�IǌӾ?�;c�"��=�@g�R#?�N�c���#���t�ߘ�qkx?"��C*���RuNQ                                                                                                                                                �`9zE[�����������[~S�²�B:U/�{��8/7(�=���{�q�<�b�e9�>.��%	���<��Z�����gM|�,��N>V��NS��fl���)�W�Z�>�c���1=T�>1�5���Njg[>x����                                                                                                                                                ?�R���ȾN-�&!|����?���(�G,���f_'�Ҿ����ǥ1�㲝Z��<�u����>j�bȢr��O�dq-� �=��c�
��>��X���"��m~|>�:?��ȾzN�X/?�",z���
/D��!��x��0���\T>���Կ���Ș�?���j�u��0����(?@�х:�@�1o�  >�%f;�� >��$�����	{�`�D�{ �g޿S/�LX��	�"}�fB���ঝ觿�P���@���o������.�U<Ɗ�                                                                                                                                                                                                                                                                                                ?�&Q�@  >�Wa~�� >�5�������t���= �1�UiLI���	���w̿���1�~y��P�jA�@������N�(�.�y^�@�>���?����~��H�"�+h�@��[iʡ>�pQ���|��Ó�g�A`!F��?�C�PXIZ� ���7��с�&�vA!�d�OG�(����:N?�'\�>x�?F9Mтee����!u�&?R��r\d�	� RĵܿF�h��0��u�spQ�?�^��+�?���9-S�@��AV�<�ۯ�4ݐm@F�jު@B�.���>�^O�S���Ҟ߰�al@����C��
o�N0�6�C3q��������B�ڿ�rS`�?��{�r���Uȿ�A
��<�9@(� ��%@]b����=��y>Q�              @�K��+>��3�xJR@���	| f@��8�%wA��xt   @�8`uR�N@�����d@V|�����@#�q��_>+��?�ޠ?���$/u�]b�    ?��g��  B�a̋H�@����M+�'�0��^��(�ޔcg���+2^W��|���p?���\�ҧ        =`L&D#�h?hj�N�M?B+R?�a߽��f I����g ������?M��֩=����^X=�gh>�'�?�N���G�@<�%��	@�\Il�V�@#�q���>/�MY�?���$/u?�ޠ?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�k���5]@�o��o? 	�a7<@�ۨjz@?�K6n�V@���_                                                =�����e�@��!8h�?����C��t[�[I�>UHJ��?TQz J�=����WL�?��i٤??@!{"���F�m�oB�=���H�?�5�ʽ��z��?��[����5����><f��^]�>r?��,m��G�(0                                                                                                                                                <�m,�X�><��<{�=�s	�s��3Ɔ��<rb��G=p�_�:G</�X�5,�>6�4�1L=���Pi�4���[Wܒ�<kpm}�A�=� ���u]<3�fBQ\�="�� ��>��T�p��� [)3��1%�ȓ>wɁ���7                                                                                                                                                �D���OM>�9�[���b�xXީl���۾��	���>e�p�%���D�j3T>�_���o>2JW{�P�>w�oxԭ���ߍb>�E*M8�+�{�l>39oԽ�	I��$���5��Լ�|��<g'>`�S����+�kjs�>3#�
�C=�
)�v�>��ڞ^�+�҆�>1�p�@&\*Y�� >7�M��  ��▲Ū���ҫ�Z5�������ڠ3���@m��  >F�F�_@ ?T7�'?���A���M��]+�[)���                                                                                                                                                                                                                                                                                                ��IQ�  >H���q  �����i����b����?o�X6��Sk�<$��)�C�  >Qܢ`  ?T$�m?���qt���M�7�ƿ[#giR�@Bsr�gu�R�jE?[�>�O�@��@o�>�w�d�i�>ٸ�?E��@Hťޭ�(�`����U~�d�>w
�� ��f�xA)M�I��I?t�w�ͷ���'4٦>8��F�=�N�<c�[\�J<��?o	� <�g9Z5tӾ��.:��:>B�u����2���8w�?�����$���$#���z�]C��:���dFc��w=z$MM��=�?,UŅ?� "�k���C�-��T��SR���#�)J�8�>Ft�)j�?T��"�?����%�@I�Ο�C>[gtagqBo���2>=
��� �m              @�e�����O++F2@���	| f@��8�%wA��xt   @�8`uR�NA�MІ�@V|�����@#L��{�
���fML8�?�C��~�@DB�;�aBo;шPx	�J�%G���E�8@GB�ļ�#*<^	���=w��rD���y7Dr��_e�0CPv%ca��?���3�_U        =)��5��>:����U�?L�lk��N=s�:Ý\c�#��-��7|'-t
�>�4d���Vӷ�O�=����7�>�G�rƖ�B�
�m�?����Kb�@#L��{�I���fM���@DB�;�a?�C��~�?�      @/��[W>�                                A�e��@  BL+��  BL��                           �H"J�`���4�=���K�'�ვ)NAqYM�1���N"@ӽ�AklHKz%�                                                ��l�1l��Q��<C�8.k�UȾ�FʔQ�>�X	�O?�?���j:�;���2��?�	LM#c�C�%� �>7�A�Lt%?H^{��+�?�C� '>�A4:�@?�M�M����~�Xu*>��$���<�2p�3�_B�����                                                                                                                                                �p�θ}ʽ�c^0�A�T���n��֩a�><�Y�ڪ�!=�8<��bH�)#���>(��̂�@����AJ9'<��X4��=�����>!�P�j��ٸ�:�d�$�Ru>��X{̽s�J���=�q�5�I�>r��v�*                                                                                                                                                ?�#�:nȾ�Ay��ξ��?0�-"?Hh��7����K����S>ʲ�pe�?���=� �&Z.�����Q���e�A���?�� 5�� �&�e��|�7%�˿!{��>���jr?���j�I&����(R?��T�!{��1��!�pG�/�U\�x?)AP���?�P�?�>�3�Gr$�?˩����@�B�  >���M`  ?W`-�v��F�D����]�S�k�S�!�
�
F�w����Z�@	����T@ғ�2�K��	R���q@@����h                                                                                                                                                                                                                                                                                                ?�j	̀  �#�!2�� ?W�NJ���Fwa����W�&�X?���P��
Gf�딬��0��H�@@	j�s�@ғ��v	n�	S+7m�E@@�-��@�h�O���cDn.�#�?پA�.@�*qq��@�i	F� ��|&��q�Alǫ'�W�)J���F�Yg�����)�&zA�CBO��I�G�kQ���|
J=?���*O�P�Fj��]�}ʝ�@	P� V��D�?�xG�9���-/"@�@E�d�@2p���@�q� iJ��UMM�@ez��}L@:<�@�M?	̛�*�kr,�	O)@���"(�@?񪭹Rs¿���+@��ވ�Ĭ?��9x�`��D�N8���ِK��LA��6A�D�Bk�B�o~@D͛��-=v��v�!?              @�_h-�7>���ߐ��@���	| f@��8�%wA��xt   @�8`uR�N@�$�h�\@V|�����@#H��>>�5[�"?��ߞ:%?����v�@D͘    ?�h��t  B��Jlc@�������(�:�_�����;�]J��,�0#���E\>go�?���O[V=        =`L��Ш?g��	��?B���갽����D�м�*�	2G����?�B�?L�.����=�� �߹F=���Ds�{?��?�dxP@:����[@�c7�(d�@#H���>�V�E�?����v�?��ߞ:%?�      @/��[W>�                                A�e��@  BL+��  BL��                           >粻�k�R@޿�n��? �]?Y��@�J���9M?�� k~r@�B�pE�                                                =����_��@� [e1?�s�g��[���f�>U�9M�?TD��߅/=��:�ƍ�?�n��dM?@T֭(ɽH<��%2�=�W���L?Ch ����'��D�?ŵ���O��5؄t�*>=��7s�+>r�� �(�*`�^�                                                                                                                                                <���6/>䪂n#�=�#���n��'�*�<r=׆mE�=q2 �p��<0��I�&�>6�ޙ#��=�7r��1��|�n���<k�-�ڶ=�S@�<4�[�>�<�{�݌�>����!W����T<
~��k�x�>x�S*�                                                                                                                                                ���D��>���/�C��B���¿ݤ "Tb���"Lp@��>e�;�����;7B��>���a>2�C��>w�z;V^��п�K>)�.S*�+|����>3�[	�o��W�)�V��qdN/�g�|���>`}7qcǓ�+l��u{>3�C�`��=�\����>�V}c��+�e��>2f��0�@&\*�&� >8PՕW  ����������ӈ�c0��TC��&���5j����@N��  >H�� ?T=�w��?�cq�����[-Dn��                                                                                                                                                                                                                                                                                                �<��2  >I<��� ����
�O���팈3����������8Y*{�(Қ��  >R�1�@ ?T=w�k�?�E#��\����['h��@B
/�n܋�SL4��G>��@���B@����.E�>�����%>�N|I�p�@H�J{_�af��_��d<�������5��DA(�a�}�?tҝOYN,��.M`>8���cE�=�i���Jc�\�W�2����?J<����)�޾�������>Cx����:�3�g^A�?��z�����AEH�]>	,Կd��m��=|,y��7=���N�m�?�i��E���+������&D��*i�QX��>G�p��?T<����?��)k'�@h�597�>\جj4kSB�j��=p,R�R�X              @��cr����y��K@���	| f@��8�%wA��xt   @�8`uR�N@��� �j@V|�����@#��O�	X�R���/�?��j+� @)l�����B�@�� ���Q��.De��-4ISC!�4��j��jh$W�uCF�Ub�ZI��_뛼¦��?���3�k�        =�ؽ�g�>������?L�#�h���a�qDs��u�Xݸ¾nL�P�v�>�5��=j�����S=�	k-?�m���?�7�0�?�`R�o�@#��O�G�S 3�\}@)l�����?��j+� ?�      @/��[W>�                                A�e��@  BL+��  BL��                           ��ĉO�!�N�ji�?ʅ�S���Ah"��.A?�������A]݇�HN�                                                ��� �����g�p����D��>Ɍs!���Ū+��:t?�p���>)ʏ�H�?�_)E3�?Wuf䶕=��i��>d��6ؓ�?(�|�B��=��J�U��?���"�26z"j�>�N���Gk>����߽�	Bfk�d�                                                                                                                                                ��������!ȇ������8��M<7�5ʄ���anJs=Լk����<���#I�>;þC�{=�y�j�
<-ѱv8�B<��_ȝN=�:��i�a n��1�����>�$L�����(Dȣ������`�a>���L��                                                                                                                                                @�ri1�1F���>$��F<�0?���(���w�S��^�խsU�?�U�MRm����h�����{DɗEL?a{ 0?³�U`>��-��r�0^��v�>���#�˯>#�'�׬��������ȿzY���x�>��E����,;��>�a'�1�>V���?2������,xv�����tA;U�h@$�?&�  >��m�x >˨��y����d~�aPܿ\�Xp����Ee[����Y��X�`?n�?b�?�F�F.�@��*\`}@�j�8?�/<�j<                                                                                                                                                                                                                                                                                                ?Ѥ̀  >�˶��� >˲�����cЀ6�!�Ƀ�J�"�Ep�|GR6��Z��ҋ�?n��B�
?�D~�j@��*�D���6��V�?�/<�O�d@x޳$�=c?4Q�U��տ!��S�@�����Y�"* B_K?I	 �=&�A mr�6¿��L�+�����.옢�տ�~�΄A&G|�۾�
6�5.2?�M��P`�>���/>�>X-&a���4Oą?>��ɳG
�R��.��(,�vT�_��?u����?���mz]�@����������N�?�B,s�9��1~(��(���K�ѽ>�����^@�U޷ ?���r$��BL���R���7��|B?y�\^��?�ɑ�3��@�����'@�p��7���@�ŉ;�A�QA��=m���P��              @��(�˿?I+lKt@���	| f@��8�%wA��xt   @�8`uR�N@����=�~@V|�����@#�)��T>|�_\�#�?y���@�;`=�����]��@ �������(D2G�?tB�W(��:��C�;Z���B�����0C��}�;�)B����?���3�{        =_����>��G���?L�o(o$�B�\F\����'q�}�eU�݅>�/0#)�q=��Q�o�=�Zu�NŠ? ��	rǿ��X�O(&@����%Q@#�)���>|�ѻV
@�;`=��?y���?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?�}Er+R�.3�wex��D���:AWy�W��?����os�AQ�K$��                                                >�y������1�!Ir������X���X�~Ǿ���P��?��Sz���g�!�`?�(���g?OtS~�<�=�w�l�>Ug���? 9C��l$�u����N?��c�9�R�4̇"�g>��2M>)>��`�{�
�z�t�'                                                                                                                                                <�Y���<%��t��B��Q`Q3B;������©��=�A'�J.���B0E�>7�j���!=�n�&ߔ�<_Ɏ3Y�<�_�>��=����yE<�O�f*	�2�gT���>��4�������m�.�D��K���>���#ŉ                                                                                                                                                @4�Y�r>�c5����ldWS�[?������I���5=⾶ �5Os��B���>�0�����sK�?����O�v���lO>�Z)��2�+ѥ���h���}���>Q�j��c��o�4���<:PHEB�>�$*�#�|�*�8�?���ж�HJ>K���@R>Ҹ7�u�E�*�jHf�6>���7)D@%ٕ�� >��"��  ���Mȿ���[�HOo�C9�|��q�9Ihʎ�����T��@?T+H�K�?�-�b�^@�:���!�s9ƫ�?�
��                                                                                                                                                                                                                                                                                                ?ҤR?   >��d��@ ���F��yV��W�u�����R�.w�ο9?!Ag�����T ���?T�!p�?�-�KH��@�G��B�sz7SϹ?�
V��
@y��}mR?0#�=4�����l@�#?�D�w��
�?%f��@��q�ֿj��¿�H�_����A'�gj�C��.L��:*?u��K"�>�ےy�`�Y�w����?F�����]1��p<�n~/Q5�C������?Hc�n\e?a�q���@�)�c1���0Y��?�NZ*�@.X��q��>�A��� �>� �ҟ��@g-�����ă'}���8�T̜ ���Ţ�;'�?cQ��r?��aF�@�=�Q:)�@��)���VovB���@Q)D Z��=�����|              @��YΪ~>����5@���	| f@��8�%wA��xt   @�8`uR�N@��(<z!@V|�����@#�$��>����?�uÈ:�?�ؖ_b��@Q)D    �k扣@  B�f���v@�>Qk ��)�i~e�n��h�R;7���c��������1ц|?���I��	        =_���ַ?e�f��r?C�UL����8�D1���tO�E�%���
2�?LB�L��=��a~v2=�6̒??����=@8�}E�B@�c��'9b@#�$�U>�� L�?�ؖ_b��?�uÈ:�?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�F�ј�@�'?U)7o?!8ϻ@���d���?r�-B?�@��{�u�G                                                =��a63�@e��,�i?�ʬ�ӾB�֗���,>U�+f�H]?T�k��H�=��*�s��?�7q&%�[?@��[� ֽI݇H��=���W9�<?�4��߽�3�$v��?�j��|���5���3�>?Hg���>s��a(��i����Y                                                                                                                                                <��#Ҷ>�!��	=�*1�s\��*lbLul<rz�wTx=qn%�&<1>�3���>6]սo��=�Y�z����}�<l�pE*-=����	<5z��� �<dk��g >�����b���#b�~��I�F�>xh��N�Q                                                                                                                                                �kcŷm�>B0�������̯��܎���Ͼ��s4VOz>e�Ϭ�[��j��$8�>@���>1�*kD2 >xp!����;�e�=�>֪�Sp��*c�̪�>4���ȺZ���ֿ���G���}oNpUV'>`�)V8#V�*c�T�T>4����=�|�GE>�9�ˉ�*co��>2�Qp��@&\*�� >8�)�"� ��ذ��P���m����U�����R���� �@�=�  >I{g�@ ?T�Ilz�Q?�@)��V�#�q��<�Z����                                                                                                                                                                                                                                                                                                �z�i>  >I�,�z� ��ݫF�D��n�}��X����Ծ۝l����(�;� >Sv�`  ?T�N�I?�@)�5���$tlt8�Z���F��@A����6�S�w�� >���P "@�p�#@Qm>Ǉ��|>>��+4�@H��^�#h�bZ��4�~�d�\[QX�@L�Y�A($����?t϶�fR��pwM��>97bϽ#=͹��l���^d�R꽾��~wX<Ӂ����˙~��>�>D\V��hž4��3�m?�@+�B3������a�]E�ऎ�eS`~~�|=ʭ�8 b=������?�((�ǽ����՛���۝OQ�r[�+��ڦ>J�β�k?T�*�X.�?�@
k�t@�����>_ݓ;{B2ͪ�<��=D�r�|D              @�ʪn��������V@���	| f@��8�%wA��xt   @�8`uR�N@����K@V|�����@#�j��� ��y���?���F�Y�@-����B#�� ��B0׏;�D�l[w���^��euݽĂ���KDT�H�"�d�9��WL3C�W���?���3�,�        =`��?}�>�o���\?L�:6U�=n��-�焼��Y!
��h��qm�>�Od�!끽�m�}�=���04�?�T��>"?��+���?���@/jr@#�j� ��n���@-����?���F�Y�?�      @/��[W>�                                A�e��@  BL+��  BL��                           ��P����]�ҷ2�_@�V�Y���Ap�n��?��Q@"QPAa	V`��                                                �R����m�vY��臿��P�����}j��(f?'�5Ro��?��-��ɶ>��8�d�?��P���S?c֢X��6����B�Q-?�q�8��?a���>�Z!��?�?M�J��1IV+�|n>�[��j�o>���[�T�1ɳ�I                                                                                                                                                �o�XjU�-�b�>���u�	�'���;v��=D��ih=�(��*?=o�m�&('>@�a�5��=���λ���%£�_d=�{ɻnV�=�Hl�F���3��1e����>��i��Ƚ"��O� �[�9!W�>�	_"��                                                                                                                                                @!D
F�8�b(~�9j���.�/�?��n���H���}�� ?7U�Â@s�@��d-��'��~w9��m�j�N����@�.3��\�ekh���3�՗ʂ�?b_���vJ���q�Կɉ1�!�?�Z�7Ύ$�,�䊇�?�Gw��?:�j;��,?���^���,�P��?����i�N@$E��  >�z�)�  ?vT������� �(4�b�r��>�H���R����m�,��HG�9Jd?��+�V�@���t���ӽ��̿�@���'�                                                                                                                                                                                                                                                                                                ?��y��  ��c�ʈ  ?u�F=] �����*���YJ{���?����u���C�3|��[�
X?������@��5[�����/-���!��%�O@��m}!�d(Hf*��@���@���奤>@��EBJ��d>��u�;A��=<�%�N���W�*��%�qb��s�ޘ�HA%-sĻߞ�a��44��ݥm�?�;X�=�w�ՋK�^����/��S��.m��0?�^'"�Y���
	W?��6|������y��@��ֈ�fS���D������]�� ��IӍK`��?�UK����j-��Q,�@��nP��}��1f�}o?�}e!�{� �zXL�x��a�3}�?��Oճ�@�x��U��@��@����?�ŕ�>SA��h)��= (pL���              @��k�:>�\�"K"�@���	| f@��8�%wA��xt   @�8`uR�N@�Ndi{�@V|�����@#�|^>3�=�c�5��?s�3���@R��q��A��
��  A9S�Ö�5D#@�J�B�#�����.[-4�G W���C�*j~�)BZ�3�_��?���3�8�        =!x3:��>�c�TQs?L��TB:ԽNQz��N�����ݹy��M9BFi>���1��G=�Á�h~T=�J�Z�2�?&��XU���g:(Ӟ�?�l��<@#�|^>4>=�d�|�@R��q��?s�3���?�      @/��[W>�                                A�e��@  BL+��  BL��                           ?�U�2��'�t��@�?W��c ٕAP_5�l?��s��fAJ���	Wc                                                >� Gr�.��+�(߿�+z�$���eNJr�Ӿ��R∭?�߻$�J=�=~-.�?�}����N?M"ѭhMýU;+��y�>Mߕ�m�?@-B�7ؽ�.�80�?��h���4{|z�Di>��P���>�Ɣ���%�
Ϫɣ�                                                                                                                                                <�:�Q�q$��=��K�{0F��z�F[��pp���=�sW��.<5P'�>6���\W=������L�˔�f�^<�g��q�I=�L�P���<r�M�/�2򚨛��>�&������G~YϽBi
�O^>��a�XO                                                                                                                                                ?�ҕ��S�>��~��ɾu7/��?��̕��o����벮���R[|M��;���>n���" �����7�f>?�c�Zt��ߧ<��L����h�*z�o�d�>"�Ow
��%ӔӀ��H�,V-/2rG>����Y��)��\X/�>!3l��r�>B�v��dW>��Ǖ �O�)��lK�ξD0��~@&3ˀ >��V��� �pg 'lH.���yv�j�5��cW[ �2І'����?>�٠?3BK�W0?��{���@�fG�;��."��_����]���I                                                                                                                                                                                                                                                                                                ?�X��  >����u`����@Ⱥ����?/T���׌���(�2���r]��F�2�@?3CHTЮ�?���  CJ@�fb0�� �.b׷֢���^n{{;@����7�?ċ�U�_�� R��(@�f�}����-M������Wc"`@�s���C-�L������EZG��c��}�A'7O�#�?��ilŻ?����&�>�^,�d�ʾsJk?	��?m�[r����q�T�w,TS>���'owUϞ?38���L�?4J5�@�@�q�����$�M{�?�kKK!��@>`+��o>�܀)|@u���JHY�@[{~��y����g��Q�3��2���؝ZRf�?B��*�R�?��� Q�@�3��/@�L�%%?Y��n�m@E�[	�v�=u��L�M�              @�	��K�>�V�1@���	| f@��8�%wA��xt   @�8`uR�N@�������@V|�����@#����*>y����\?�0��;?�Uǹw�@E�X    ?��X�  B�8��^�@�F^�C��*ϔL-;8������)�ҴX������Sϓ�a?���'>�0        =_T�bͅ?dZ�M�}�?C�����y����΋�.��f|��ۿv"P�?K�5V��'=��#���!=�Q�c��J?/J��@6Ӌ�DH@�\�O��@#�����>y��O��?�Uǹw�?�0��;?�      @/��[W>�                                A�e��@  BL+��  BL��                           >���ܯ�@ߙ��`l?^����@��X~?
r	��@��f̝<                                                =����=@1?�_?�.q�Y��=�Zz��>VިQu?T�b�tK�=���qЃ5?�R�ͅ�?@�䞸�K��e�&=��m�Z?���t�N��ِ�V�?�%�O0�5�߇N�>@t%���>twR&������?9�                                                                                                                                                <���� �>+�~��=����OY��h$�<r��mK=q�ϱ��<1����d>6mffM=��9������r��(<l}�����=�#pS�A<6V=�����<�	V[�>��}�1༵ϸ��X���!vHS!`>x�h%8cp                                                                                                                                                ��]���>���ٽ���ݿۑ�� ۾�4w��W�>e�������V.�>6�5��>1���yC�>xy:�nk����R��>�!���x�)������>4�R�&(��%�������KC�پ~LA���>`��)��)��5�i>4�7Um�W=��<dv>h)0l�2�)ǟ�t��>3��$EO�@&\+37� >9�<��  ���KD>A��<۾��Ҿ����#}�ܧ���@�4�&  >K�<E� ?Tδ4���?����w��@�1a�[ ��L��                                                                                                                                                                                                                                                                                                ��%�  >J�x�� ���Ze�����=�����2>�
ԕ��ZQ��R�(�F�� >Tm�A� ?Tθ��?�� ��q�����Q��[ �e�RI@A0�����T`=;?ڂ>��K��6,@�?��U	�>�4�E�p>ۿb��*�@H��<�7ƾcdZ2���d�m��w���M�\`A'��$@?t�������MM�
h>9����b�=��6�5�`1�&�.G��2?
M��<�9���`Z�Σ|"|��>ER��/U�6<p�bm1?����� ��lB�Q��]Y�چ�n�e�8X{f=�����<=�6q�T�h?��킏ƾ�7�)`쀾�Z1n����-J��نo>Lpp��G?TΒW??�t�^A@I`�~A%>`Đ� @,}��]=Z@����6              @�c��]ac>��	6���@���	| f@��8�%wA��xt   @�8`uR�N@�w!YN��@V|�����@$ `=di�> �ã�
?��еg?���0�Ʊ�,}�    ?�J��X  B�ǡ��/�@�9ო*�,H�Yv�N��l�_rv����ɠ��'����?�����        =^���bΝ?b���>?D%�Yt��6D�������w9־ڕ����]?J�%^� _=��3��=����wL"?}��J�@4���I��@�JD�Ǝ@$ `=dam> �3!'1?���0�Ʊ?��еg?�      @/��[W>�                                A�e��@  BL+��  BL��                           >�I����@��z�T�?�d��@�`��f�?'_��@�z�w4                                                =�i?�?@ �y����?ʋ#�������:1*>V|��?UY#�=����{?��5�W�?@��^�G�M��SI�=�R8Qq �?ۤ�������"a��?����j�5բ�n;>Aia�G�U>ui!wj����s���                                                                                                                                                <�G�
�>�~z=��pӻ�`�t��`<sz0g��=q揤|�<2���r>5���J(=�Y�@����-A�Ŀ�<l��:�_=�gt>�<7Y)���6�;��e;��>���������:i��b�"��>y0��PG                                                                                                                                                ������>��.C ��m���> �ڌpF��ᾤ�=�ą>e�f��Q��:�ܨU>�y1\��>1�P_�%N>y	�apTH�k�R/5�>t��B��)%n�R>5Y�-���ɪV�Vῴ�y2)�e�<�DY>`��ra8�)$���e�>5YgC~Q�=�%[֌6>օN���)$�il�>48�=��k@&\+W�� >:e@ƀ ��p�S�-��	6|fü��	%l�<�݈�QD@2|�  >L�1)�@ ?U.���?��ҍrL� +��|��[�� ��                                                                                                                                                                                                                                                                                                �(�A�  >K}$��� ����31��
3��k������4���;��_=��(�m�À >U����  ?U.���F�?��7?7� j<֡��[�4��g@@Åp�NܾU�-nH�>�$��:��@��R
>��v;=2>ܠ	P��@H�͸�~�d����[�e.5�H���=A' op);-?t����~>��w/>:��a���=�S��C��ak�ž����O��<ܴ��ԧ��Kz����>F�3�p�ؾ8$�4Of?��:--��,Q��J�]����ƿf�c1�w=��tO�X=�Ll%��?�(�b�O򾯢uЩI־�;������/�Yyō>O�����?U.Y���a?��q�Xߩ@5?]�>bQ��.��    ��           PLASMA        4     h  h                                            	                                                      4  �                  DENE   DENI   BMAG   SPECIES    LABEL      LABELS        P  �                                                  `                                            	          	                                                 (          0          8          @          H          NAME   AMU    ZCHARGE    FRAC   TEMPPAR    AA     BB     DD     VD     A$@WVA$@WVG:5       H+  ?�      ?�      ?�z�0�?��@   ?�      ?�      ?�                    O+  @/��`   ?�      ?�\(�x�w?��@   ?�      ?�      ?�                    e-  ?Aد��f��      ?�      ?*6��   ?�      ?�      ?�                    e+          ?�              ?�      ?�      ?����   ?�                    e+          ?�              ?�      ?�      ?����   ?�                    e+          ?�              ?�      ?�      ?����   ?�                 G   GDENe=2.47e+05cm!u-3!n B!d0!n=4.77e+04 nT  0.0200 H+, 0.980 O+, 1.00 e-,    9   90.0200 H+ T=9.00e-05 keV A=1.00 B=0.500 D=1.00 V=0.00 m/s      8   80.980 O+ T=9.00e-05 keV A=1.00 B=0.500 D=1.00 V=0.00 m/s   7   71.00 e- T=0.000200 keV A=1.00 B=0.500 D=1.00 V=0.00 m/s    3   30.00 e+ T=1.00 keV A=1.00 B=0.100 D=1.00 V=0.00 m/s    3   30.00 e+ T=1.00 keV A=1.00 B=0.100 D=1.00 V=0.00 m/s    3   30.00 e+ T=1.00 keV A=1.00 B=0.100 D=1.00 V=0.00 m/s                